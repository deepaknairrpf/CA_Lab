module main_memory (en,w, addr, dataIn, dataOut, clk);





input w,en,clk;
input [31:0]dataIn;
input [11:0]addr;
output reg [127:0] dataOut;


reg [32:0]memory[4095:0];
wire [11:0] w1,w2,w3,w4;




assign w1[11:2] = addr[11:2];
assign w2[11:2] = addr[11:2];
assign w3[11:2] = addr[11:2];
assign w4[11:2] = addr[11:2];

assign w1[1:0] = 2'b00;
assign w2[1:0] = 2'b01;
assign w3[1:0] = 2'b10;
assign w4[1:0] = 2'b11;






always@(negedge clk)
begin

if (en==1)
begin

    if (w==1)
        memory[addr] <= dataIn;
        
    else
    begin
    
        dataOut[127:96] <= memory[w1];
        dataOut[95 :64] <= memory[w2];
        dataOut[63 :32] <= memory[w3];
        dataOut[31 :0 ] <= memory[w4];
        
        
    end  

end
end


initial
begin

memory[0] = 32'd4289383;
memory[1] = 32'd6930886;
memory[2] = 32'd1692777;
memory[3] = 32'd4636915;
memory[4] = 32'd7747793;
memory[5] = 32'd4238335;
memory[6] = 32'd9885386;
memory[7] = 32'd9760492;
memory[8] = 32'd6516649;
memory[9] = 32'd9641421;
memory[10] = 32'd5202362;
memory[11] = 32'd490027;
memory[12] = 32'd3368690;
memory[13] = 32'd2520059;
memory[14] = 32'd4897763;
memory[15] = 32'd7513926;
memory[16] = 32'd5180540;
memory[17] = 32'd383426;
memory[18] = 32'd4089172;
memory[19] = 32'd3455736;
memory[20] = 32'd5005211;
memory[21] = 32'd1595368;
memory[22] = 32'd4702567;
memory[23] = 32'd6956429;
memory[24] = 32'd6465782;
memory[25] = 32'd1021530;
memory[26] = 32'd8722862;
memory[27] = 32'd3665123;
memory[28] = 32'd5174067;
memory[29] = 32'd8703135;
memory[30] = 32'd1513929;
memory[31] = 32'd1979802;
memory[32] = 32'd5634022;
memory[33] = 32'd5723058;
memory[34] = 32'd9133069;
memory[35] = 32'd5898167;
memory[36] = 32'd9961393;
memory[37] = 32'd9018456;
memory[38] = 32'd8175011;
memory[39] = 32'd6478042;
memory[40] = 32'd1176229;
memory[41] = 32'd3377373;
memory[42] = 32'd9484421;
memory[43] = 32'd4544919;
memory[44] = 32'd8413784;
memory[45] = 32'd6898537;
memory[46] = 32'd4575198;
memory[47] = 32'd3594324;
memory[48] = 32'd9798315;
memory[49] = 32'd8664370;
memory[50] = 32'd9566413;
memory[51] = 32'd4803526;
memory[52] = 32'd2776091;
memory[53] = 32'd4268980;
memory[54] = 32'd1759956;
memory[55] = 32'd9241873;
memory[56] = 32'd7806862;
memory[57] = 32'd2999170;
memory[58] = 32'd2906996;
memory[59] = 32'd5497281;
memory[60] = 32'd1702305;
memory[61] = 32'd4420925;
memory[62] = 32'd7477084;
memory[63] = 32'd7336327;
memory[64] = 32'd2660336;
memory[65] = 32'd9126505;
memory[66] = 32'd5750846;
memory[67] = 32'd2621729;
memory[68] = 32'd661313;
memory[69] = 32'd3925857;
memory[70] = 32'd1616124;
memory[71] = 32'd4353895;
memory[72] = 32'd9819582;
memory[73] = 32'd1100545;
memory[74] = 32'd8898814;
memory[75] = 32'd8233367;
memory[76] = 32'd515434;
memory[77] = 32'd5990364;
memory[78] = 32'd4344043;
memory[79] = 32'd313750;
memory[80] = 32'd7171087;
memory[81] = 32'd6426808;
memory[82] = 32'd5117276;
memory[83] = 32'd9947178;
memory[84] = 32'd695788;
memory[85] = 32'd9393584;
memory[86] = 32'd1705403;
memory[87] = 32'd8502651;
memory[88] = 32'd2392754;
memory[89] = 32'd4612399;
memory[90] = 32'd3999932;
memory[91] = 32'd4095060;
memory[92] = 32'd1549676;
memory[93] = 32'd3993368;
memory[94] = 32'd3947739;
memory[95] = 32'd4210012;
memory[96] = 32'd5636226;
memory[97] = 32'd9698586;
memory[98] = 32'd9348094;
memory[99] = 32'd6297539;
memory[100] = 32'd6140795;
memory[101] = 32'd3480570;
memory[102] = 32'd651434;
memory[103] = 32'd5960378;
memory[104] = 32'd7097467;
memory[105] = 32'd2066601;
memory[106] = 32'd6710097;
memory[107] = 32'd7612902;
memory[108] = 32'd573317;
memory[109] = 32'd3570492;
memory[110] = 32'd7926652;
memory[111] = 32'd260756;
memory[112] = 32'd9997301;
memory[113] = 32'd5560280;
memory[114] = 32'd2724286;
memory[115] = 32'd3209441;
memory[116] = 32'd4953865;
memory[117] = 32'd4429689;
memory[118] = 32'd4228444;
memory[119] = 32'd7346619;
memory[120] = 32'd1558440;
memory[121] = 32'd744729;
memory[122] = 32'd3958031;
memory[123] = 32'd3108117;
memory[124] = 32'd4738097;
memory[125] = 32'd7905771;
memory[126] = 32'd9834481;
memory[127] = 32'd2890675;
memory[128] = 32'd120709;
memory[129] = 32'd1698927;
memory[130] = 32'd1704567;
memory[131] = 32'd8777856;
memory[132] = 32'd5179497;
memory[133] = 32'd4872353;
memory[134] = 32'd7254586;
memory[135] = 32'd2276965;
memory[136] = 32'd9455306;
memory[137] = 32'd3964683;
memory[138] = 32'd2406219;
memory[139] = 32'd28624;
memory[140] = 32'd51528;
memory[141] = 32'd332871;
memory[142] = 32'd2805732;
memory[143] = 32'd48829;
memory[144] = 32'd8409503;
memory[145] = 32'd5530019;
memory[146] = 32'd3258270;
memory[147] = 32'd3363368;
memory[148] = 32'd9959708;
memory[149] = 32'd7486715;
memory[150] = 32'd3226340;
memory[151] = 32'd1518149;
memory[152] = 32'd747796;
memory[153] = 32'd9700723;
memory[154] = 32'd7142618;
memory[155] = 32'd8002245;
memory[156] = 32'd122846;
memory[157] = 32'd9493451;
memory[158] = 32'd892921;
memory[159] = 32'd243555;
memory[160] = 32'd1192379;
memory[161] = 32'd2597488;
memory[162] = 32'd1537764;
memory[163] = 32'd8888228;
memory[164] = 32'd7469841;
memory[165] = 32'd8792350;
memory[166] = 32'd1165193;
memory[167] = 32'd9441500;
memory[168] = 32'd2757034;
memory[169] = 32'd6087764;
memory[170] = 32'd9470124;
memory[171] = 32'd5324914;
memory[172] = 32'd8936987;
memory[173] = 32'd2275856;
memory[174] = 32'd5373743;
memory[175] = 32'd7346491;
memory[176] = 32'd322227;
memory[177] = 32'd1148365;
memory[178] = 32'd709859;
memory[179] = 32'd281936;
memory[180] = 32'd1151432;
memory[181] = 32'd6452551;
memory[182] = 32'd4316437;
memory[183] = 32'd1899228;
memory[184] = 32'd6153275;
memory[185] = 32'd3975407;
memory[186] = 32'd9901474;
memory[187] = 32'd6276121;
memory[188] = 32'd3468858;
memory[189] = 32'd794395;
memory[190] = 32'd9036029;
memory[191] = 32'd4661237;
memory[192] = 32'd5908235;
memory[193] = 32'd573793;
memory[194] = 32'd6065818;
memory[195] = 32'd5894428;
memory[196] = 32'd9366143;
memory[197] = 32'd7231011;
memory[198] = 32'd5335928;
memory[199] = 32'd4639529;
memory[200] = 32'd3318776;
memory[201] = 32'd7322404;
memory[202] = 32'd9964443;
memory[203] = 32'd2255763;
memory[204] = 32'd2114613;
memory[205] = 32'd7854538;
memory[206] = 32'd2118606;
memory[207] = 32'd2436840;
memory[208] = 32'd9002904;
memory[209] = 32'd5344818;
memory[210] = 32'd5235128;
memory[211] = 32'd2670688;
memory[212] = 32'd1797369;
memory[213] = 32'd2067917;
memory[214] = 32'd4569917;
memory[215] = 32'd466996;
memory[216] = 32'd6043324;
memory[217] = 32'd6987743;
memory[218] = 32'd9259470;
memory[219] = 32'd9512183;
memory[220] = 32'd298490;
memory[221] = 32'd8295499;
memory[222] = 32'd6689772;
memory[223] = 32'd6206725;
memory[224] = 32'd1385644;
memory[225] = 32'd2755590;
memory[226] = 32'd4617505;
memory[227] = 32'd3268139;
memory[228] = 32'd2502954;
memory[229] = 32'd2469786;
memory[230] = 32'd7907669;
memory[231] = 32'd8338082;
memory[232] = 32'd2308542;
memory[233] = 32'd388464;
memory[234] = 32'd3110197;
memory[235] = 32'd6939507;
memory[236] = 32'd759355;
memory[237] = 32'd5228804;
memory[238] = 32'd9376348;
memory[239] = 32'd2278611;
memory[240] = 32'd573622;
memory[241] = 32'd7127828;
memory[242] = 32'd4949299;
memory[243] = 32'd4887343;
memory[244] = 32'd9195746;
memory[245] = 32'd2035568;
memory[246] = 32'd5354340;
memory[247] = 32'd7755422;
memory[248] = 32'd9023311;
memory[249] = 32'd4613810;
memory[250] = 32'd7267605;
memory[251] = 32'd9321801;
memory[252] = 32'd5425661;
memory[253] = 32'd6473730;
memory[254] = 32'd8044878;
memory[255] = 32'd6811305;
memory[256] = 32'd9229320;
memory[257] = 32'd5178736;
memory[258] = 32'd79444;
memory[259] = 32'd4248626;
memory[260] = 32'd7648522;
memory[261] = 32'd503465;
memory[262] = 32'd2586708;
memory[263] = 32'd2473416;
memory[264] = 32'd3408282;
memory[265] = 32'd8213258;
memory[266] = 32'd9412924;
memory[267] = 32'd4167637;
memory[268] = 32'd3442062;
memory[269] = 32'd1305624;
memory[270] = 32'd8962600;
memory[271] = 32'd6532036;
memory[272] = 32'd8433452;
memory[273] = 32'd3911899;
memory[274] = 32'd1419379;
memory[275] = 32'd145550;
memory[276] = 32'd5947468;
memory[277] = 32'd9290071;
memory[278] = 32'd7900973;
memory[279] = 32'd7487131;
memory[280] = 32'd3903881;
memory[281] = 32'd7684930;
memory[282] = 32'd6808933;
memory[283] = 32'd1845894;
memory[284] = 32'd4158660;
memory[285] = 32'd7370163;
memory[286] = 32'd8657199;
memory[287] = 32'd3387981;
memory[288] = 32'd2548899;
memory[289] = 32'd1252996;
memory[290] = 32'd152959;
memory[291] = 32'd2713773;
memory[292] = 32'd4272813;
memory[293] = 32'd2739668;
memory[294] = 32'd5187190;
memory[295] = 32'd7681095;
memory[296] = 32'd952926;
memory[297] = 32'd7116466;
memory[298] = 32'd4365084;
memory[299] = 32'd6911340;
memory[300] = 32'd8422090;
memory[301] = 32'd3327684;
memory[302] = 32'd3443376;
memory[303] = 32'd6855542;
memory[304] = 32'd9755936;
memory[305] = 32'd7379107;
memory[306] = 32'd9517445;
memory[307] = 32'd8219756;
memory[308] = 32'd6669179;
memory[309] = 32'd7418418;
memory[310] = 32'd5706887;
memory[311] = 32'd3089412;
memory[312] = 32'd5103348;
memory[313] = 32'd5032172;
memory[314] = 32'd7451659;
memory[315] = 32'd9262009;
memory[316] = 32'd2402336;
memory[317] = 32'd8625210;
memory[318] = 32'd5166342;
memory[319] = 32'd7467587;
memory[320] = 32'd9878206;
memory[321] = 32'd5319301;
memory[322] = 32'd2697713;
memory[323] = 32'd6667372;
memory[324] = 32'd575321;
memory[325] = 32'd401255;
memory[326] = 32'd6864819;
memory[327] = 32'd4044599;
memory[328] = 32'd7517721;
memory[329] = 32'd1229904;
memory[330] = 32'd955939;
memory[331] = 32'd5939811;
memory[332] = 32'd7073940;
memory[333] = 32'd6915667;
memory[334] = 32'd5311705;
memory[335] = 32'd9346228;
memory[336] = 32'd6811127;
memory[337] = 32'd4829150;
memory[338] = 32'd7565984;
memory[339] = 32'd5996658;
memory[340] = 32'd4763920;
memory[341] = 32'd5789224;
memory[342] = 32'd1602422;
memory[343] = 32'd9867269;
memory[344] = 32'd821396;
memory[345] = 32'd9054081;
memory[346] = 32'd1645630;
memory[347] = 32'd5740084;
memory[348] = 32'd7679292;
memory[349] = 32'd6811972;
memory[350] = 32'd3207672;
memory[351] = 32'd73850;
memory[352] = 32'd4647625;
memory[353] = 32'd5905385;
memory[354] = 32'd6741222;
memory[355] = 32'd7739299;
memory[356] = 32'd6306640;
memory[357] = 32'd3606042;
memory[358] = 32'd1783898;
memory[359] = 32'd6340713;
memory[360] = 32'd7352298;
memory[361] = 32'd5256190;
memory[362] = 32'd2280524;
memory[363] = 32'd6942590;
memory[364] = 32'd4688209;
memory[365] = 32'd108581;
memory[366] = 32'd6288819;
memory[367] = 32'd1499336;
memory[368] = 32'd4937732;
memory[369] = 32'd6371155;
memory[370] = 32'd7495994;
memory[371] = 32'd2218004;
memory[372] = 32'd2160379;
memory[373] = 32'd1614769;
memory[374] = 32'd2085273;
memory[375] = 32'd2981776;
memory[376] = 32'd668850;
memory[377] = 32'd6247255;
memory[378] = 32'd8721860;
memory[379] = 32'd8348142;
memory[380] = 32'd5575579;
memory[381] = 32'd4445884;
memory[382] = 32'd8421993;
memory[383] = 32'd223205;
memory[384] = 32'd2867621;
memory[385] = 32'd7679567;
memory[386] = 32'd7962504;
memory[387] = 32'd1690613;
memory[388] = 32'd3801961;
memory[389] = 32'd2262754;
memory[390] = 32'd8031326;
memory[391] = 32'd1154259;
memory[392] = 32'd7518944;
memory[393] = 32'd2828202;
memory[394] = 32'd613202;
memory[395] = 32'd4723506;
memory[396] = 32'd2936784;
memory[397] = 32'd6902021;
memory[398] = 32'd6222842;
memory[399] = 32'd390868;
memory[400] = 32'd5789528;
memory[401] = 32'd6235189;
memory[402] = 32'd2608872;
memory[403] = 32'd7949908;
memory[404] = 32'd7849958;
memory[405] = 32'd7210498;
memory[406] = 32'd3448036;
memory[407] = 32'd8518808;
memory[408] = 32'd3457753;
memory[409] = 32'd4686248;
memory[410] = 32'd9383303;
memory[411] = 32'd9033333;
memory[412] = 32'd9132133;
memory[413] = 32'd321648;
memory[414] = 32'd1772890;
memory[415] = 32'd1999754;
memory[416] = 32'd517567;
memory[417] = 32'd2251746;
memory[418] = 32'd3690368;
memory[419] = 32'd4319529;
memory[420] = 32'd4514500;
memory[421] = 32'd4238046;
memory[422] = 32'd5473788;
memory[423] = 32'd4549797;
memory[424] = 32'd7066249;
memory[425] = 32'd6086990;
memory[426] = 32'd9273303;
memory[427] = 32'd3033;
memory[428] = 32'd5505363;
memory[429] = 32'd8012497;
memory[430] = 32'd2910253;
memory[431] = 32'd1294892;
memory[432] = 32'd4247686;
memory[433] = 32'd5519125;
memory[434] = 32'd1761152;
memory[435] = 32'd4613996;
memory[436] = 32'd5245975;
memory[437] = 32'd5209188;
memory[438] = 32'd5649157;
memory[439] = 32'd8703729;
memory[440] = 32'd9895436;
memory[441] = 32'd5032460;
memory[442] = 32'd253414;
memory[443] = 32'd1543921;
memory[444] = 32'd7870460;
memory[445] = 32'd2026304;
memory[446] = 32'd6060028;
memory[447] = 32'd8388027;
memory[448] = 32'd4278050;
memory[449] = 32'd2266748;
memory[450] = 32'd2707556;
memory[451] = 32'd1308902;
memory[452] = 32'd6504794;
memory[453] = 32'd697697;
memory[454] = 32'd5858699;
memory[455] = 32'd3571043;
memory[456] = 32'd9301039;
memory[457] = 32'd5132002;
memory[458] = 32'd6090428;
memory[459] = 32'd4806403;
memory[460] = 32'd3144500;
memory[461] = 32'd9000681;
memory[462] = 32'd8617647;
memory[463] = 32'd9908538;
memory[464] = 32'd7036159;
memory[465] = 32'd2895151;
memory[466] = 32'd4522535;
memory[467] = 32'd2282134;
memory[468] = 32'd8104339;
memory[469] = 32'd171692;
memory[470] = 32'd3502215;
memory[471] = 32'd516127;
memory[472] = 32'd7720504;
memory[473] = 32'd3755629;
memory[474] = 32'd2060049;
memory[475] = 32'd5590964;
memory[476] = 32'd8298285;
memory[477] = 32'd636429;
memory[478] = 32'd6495343;
memory[479] = 32'd2576335;
memory[480] = 32'd2903177;
memory[481] = 32'd9202900;
memory[482] = 32'd3885238;
memory[483] = 32'd9407971;
memory[484] = 32'd2416949;
memory[485] = 32'd2260289;
memory[486] = 32'd5495367;
memory[487] = 32'd1717988;
memory[488] = 32'd7392292;
memory[489] = 32'd1585795;
memory[490] = 32'd9040743;
memory[491] = 32'd3053144;
memory[492] = 32'd3102829;
memory[493] = 32'd7658390;
memory[494] = 32'd2961682;
memory[495] = 32'd2655340;
memory[496] = 32'd553541;
memory[497] = 32'd569;
memory[498] = 32'd7453826;
memory[499] = 32'd1174232;
memory[500] = 32'd172261;
memory[501] = 32'd956042;
memory[502] = 32'd1690360;
memory[503] = 32'd409117;
memory[504] = 32'd7228023;
memory[505] = 32'd6266761;
memory[506] = 32'd6000081;
memory[507] = 32'd5526309;
memory[508] = 32'd6903190;
memory[509] = 32'd2495425;
memory[510] = 32'd618996;
memory[511] = 32'd9806367;
memory[512] = 32'd4214677;
memory[513] = 32'd4504234;
memory[514] = 32'd1730690;
memory[515] = 32'd6631626;
memory[516] = 32'd6764524;
memory[517] = 32'd7226057;
memory[518] = 32'd8349614;
memory[519] = 32'd6673168;
memory[520] = 32'd1328205;
memory[521] = 32'd7390358;
memory[522] = 32'd9726312;
memory[523] = 32'd6947386;
memory[524] = 32'd7565100;
memory[525] = 32'd5204346;
memory[526] = 32'd9602726;
memory[527] = 32'd634994;
memory[528] = 32'd5204916;
memory[529] = 32'd7056552;
memory[530] = 32'd4325578;
memory[531] = 32'd7893529;
memory[532] = 32'd528946;
memory[533] = 32'd8532290;
memory[534] = 32'd8302647;
memory[535] = 32'd7756970;
memory[536] = 32'd4799051;
memory[537] = 32'd6819080;
memory[538] = 32'd5799631;
memory[539] = 32'd4218593;
memory[540] = 32'd1830857;
memory[541] = 32'd6418627;
memory[542] = 32'd6541312;
memory[543] = 32'd8561886;
memory[544] = 32'd3439214;
memory[545] = 32'd788355;
memory[546] = 32'd5193512;
memory[547] = 32'd2720090;
memory[548] = 32'd8014412;
memory[549] = 32'd6059479;
memory[550] = 32'd1909610;
memory[551] = 32'd1858969;
memory[552] = 32'd5966189;
memory[553] = 32'd4152274;
memory[554] = 32'd8806355;
memory[555] = 32'd6047641;
memory[556] = 32'd9356620;
memory[557] = 32'd925433;
memory[558] = 32'd9198987;
memory[559] = 32'd7077888;
memory[560] = 32'd498338;
memory[561] = 32'd3524566;
memory[562] = 32'd7487770;
memory[563] = 32'd1027284;
memory[564] = 32'd2056856;
memory[565] = 32'd5790417;
memory[566] = 32'd1300606;
memory[567] = 32'd9372260;
memory[568] = 32'd5125849;
memory[569] = 32'd7100237;
memory[570] = 32'd6107205;
memory[571] = 32'd9473059;
memory[572] = 32'd6035217;
memory[573] = 32'd2648518;
memory[574] = 32'd8034945;
memory[575] = 32'd1990783;
memory[576] = 32'd3436873;
memory[577] = 32'd3228458;
memory[578] = 32'd4710873;
memory[579] = 32'd3967637;
memory[580] = 32'd1804289;
memory[581] = 32'd6620483;
memory[582] = 32'd5826607;
memory[583] = 32'd7770478;
memory[584] = 32'd772757;
memory[585] = 32'd7149314;
memory[586] = 32'd6334471;
memory[587] = 32'd2645729;
memory[588] = 32'd591100;
memory[589] = 32'd5533459;
memory[590] = 32'd9723618;
memory[591] = 32'd1089438;
memory[592] = 32'd9058025;
memory[593] = 32'd7211388;
memory[594] = 32'd4633074;
memory[595] = 32'd3631233;
memory[596] = 32'd5518157;
memory[597] = 32'd5933681;
memory[598] = 32'd3003493;
memory[599] = 32'd3160358;
memory[600] = 32'd5550270;
memory[601] = 32'd9110699;
memory[602] = 32'd2633417;
memory[603] = 32'd4101839;
memory[604] = 32'd4275569;
memory[605] = 32'd668363;
memory[606] = 32'd6092622;
memory[607] = 32'd228794;
memory[608] = 32'd6413173;
memory[609] = 32'd3319847;
memory[610] = 32'd4196431;
memory[611] = 32'd8217462;
memory[612] = 32'd2456682;
memory[613] = 32'd2539390;
memory[614] = 32'd8504292;
memory[615] = 32'd5745791;
memory[616] = 32'd2205057;
memory[617] = 32'd7355115;
memory[618] = 32'd8391521;
memory[619] = 32'd2796157;
memory[620] = 32'd2888574;
memory[621] = 32'd631491;
memory[622] = 32'd6401947;
memory[623] = 32'd4462951;
memory[624] = 32'd359231;
memory[625] = 32'd1035021;
memory[626] = 32'd610537;
memory[627] = 32'd8393740;
memory[628] = 32'd9485054;
memory[629] = 32'd3614030;
memory[630] = 32'd1554098;
memory[631] = 32'd5035325;
memory[632] = 32'd5241081;
memory[633] = 32'd4187516;
memory[634] = 32'd1653516;
memory[635] = 32'd2033002;
memory[636] = 32'd7372231;
memory[637] = 32'd7746139;
memory[638] = 32'd2261796;
memory[639] = 32'd3785404;
memory[640] = 32'd3582338;
memory[641] = 32'd8974580;
memory[642] = 32'd4519218;
memory[643] = 32'd6039021;
memory[644] = 32'd1513970;
memory[645] = 32'd5539862;
memory[646] = 32'd1784812;
memory[647] = 32'd6235379;
memory[648] = 32'd2894977;
memory[649] = 32'd2692685;
memory[650] = 32'd9031536;
memory[651] = 32'd8299904;
memory[652] = 32'd3324176;
memory[653] = 32'd5433483;
memory[654] = 32'd5279207;
memory[655] = 32'd6199759;
memory[656] = 32'd8984857;
memory[657] = 32'd5889744;
memory[658] = 32'd4593499;
memory[659] = 32'd8469911;
memory[660] = 32'd2020127;
memory[661] = 32'd8663950;
memory[662] = 32'd3505236;
memory[663] = 32'd9777560;
memory[664] = 32'd5367818;
memory[665] = 32'd7675105;
memory[666] = 32'd1810563;
memory[667] = 32'd2740049;
memory[668] = 32'd5421244;
memory[669] = 32'd6588711;
memory[670] = 32'd9041805;
memory[671] = 32'd1519934;
memory[672] = 32'd5563291;
memory[673] = 32'd6077375;
memory[674] = 32'd7558955;
memory[675] = 32'd9593614;
memory[676] = 32'd4133589;
memory[677] = 32'd9343768;
memory[678] = 32'd5828993;
memory[679] = 32'd9544918;
memory[680] = 32'd4552805;
memory[681] = 32'd7376882;
memory[682] = 32'd7844822;
memory[683] = 32'd7876982;
memory[684] = 32'd5326717;
memory[685] = 32'd3124030;
memory[686] = 32'd6593093;
memory[687] = 32'd4311574;
memory[688] = 32'd1530126;
memory[689] = 32'd1186593;
memory[690] = 32'd2781486;
memory[691] = 32'd3550253;
memory[692] = 32'd9850543;
memory[693] = 32'd8803074;
memory[694] = 32'd3327814;
memory[695] = 32'd7734713;
memory[696] = 32'd6478179;
memory[697] = 32'd5138377;
memory[698] = 32'd474762;
memory[699] = 32'd4415775;
memory[700] = 32'd1727088;
memory[701] = 32'd2032919;
memory[702] = 32'd5935710;
memory[703] = 32'd9806732;
memory[704] = 32'd8110294;
memory[705] = 32'd6011017;
memory[706] = 32'd9400346;
memory[707] = 32'd4760235;
memory[708] = 32'd7871137;
memory[709] = 32'd7745691;
memory[710] = 32'd4305153;
memory[711] = 32'd2423943;
memory[712] = 32'd5122573;
memory[713] = 32'd4666328;
memory[714] = 32'd300925;
memory[715] = 32'd449291;
memory[716] = 32'd306710;
memory[717] = 32'd6894018;
memory[718] = 32'd7277217;
memory[719] = 32'd1836836;
memory[720] = 32'd596963;
memory[721] = 32'd2575055;
memory[722] = 32'd5387090;
memory[723] = 32'd2963858;
memory[724] = 32'd1378130;
memory[725] = 32'd8714904;
memory[726] = 32'd698571;
memory[727] = 32'd372661;
memory[728] = 32'd6369633;
memory[729] = 32'd3689685;
memory[730] = 32'd7304789;
memory[731] = 32'd613073;
memory[732] = 32'd5722604;
memory[733] = 32'd5756851;
memory[734] = 32'd419805;
memory[735] = 32'd6349250;
memory[736] = 32'd1767868;
memory[737] = 32'd2336503;
memory[738] = 32'd1109485;
memory[739] = 32'd9639006;
memory[740] = 32'd82195;
memory[741] = 32'd5414639;
memory[742] = 32'd2062949;
memory[743] = 32'd7721120;
memory[744] = 32'd80967;
memory[745] = 32'd4880226;
memory[746] = 32'd686763;
memory[747] = 32'd387677;
memory[748] = 32'd4290596;
memory[749] = 32'd7963981;
memory[750] = 32'd4740865;
memory[751] = 32'd4887560;
memory[752] = 32'd539036;
memory[753] = 32'd127955;
memory[754] = 32'd367770;
memory[755] = 32'd4433518;
memory[756] = 32'd1359211;
memory[757] = 32'd1066342;
memory[758] = 32'd7322532;
memory[759] = 32'd245196;
memory[760] = 32'd7272379;
memory[761] = 32'd4627321;
memory[762] = 32'd858270;
memory[763] = 32'd2994984;
memory[764] = 32'd384172;
memory[765] = 32'd3794427;
memory[766] = 32'd9344234;
memory[767] = 32'd2152040;
memory[768] = 32'd8647283;
memory[769] = 32'd2970072;
memory[770] = 32'd4307398;
memory[771] = 32'd1245830;
memory[772] = 32'd901063;
memory[773] = 32'd6370347;
memory[774] = 32'd8966950;
memory[775] = 32'd982030;
memory[776] = 32'd1250573;
memory[777] = 32'd9653714;
memory[778] = 32'd3886059;
memory[779] = 32'd8057522;
memory[780] = 32'd134047;
memory[781] = 32'd8626924;
memory[782] = 32'd2945082;
memory[783] = 32'd3189435;
memory[784] = 32'd1271232;
memory[785] = 32'd5829204;
memory[786] = 32'd7622954;
memory[787] = 32'd2630443;
memory[788] = 32'd9411898;
memory[789] = 32'd4945486;
memory[790] = 32'd2875640;
memory[791] = 32'd6684278;
memory[792] = 32'd2089159;
memory[793] = 32'd6250262;
memory[794] = 32'd9679262;
memory[795] = 32'd4989683;
memory[796] = 32'd2561041;
memory[797] = 32'd1539848;
memory[798] = 32'd7141723;
memory[799] = 32'd1208324;
memory[800] = 32'd7026272;
memory[801] = 32'd1449122;
memory[802] = 32'd2454154;
memory[803] = 32'd7927335;
memory[804] = 32'd335821;
memory[805] = 32'd3937457;
memory[806] = 32'd8909365;
memory[807] = 32'd4102747;
memory[808] = 32'd3591171;
memory[809] = 32'd5311776;
memory[810] = 32'd2160269;
memory[811] = 32'd3725218;
memory[812] = 32'd3938701;
memory[813] = 32'd7621703;
memory[814] = 32'd6914653;
memory[815] = 32'd5209933;
memory[816] = 32'd3450907;
memory[817] = 32'd7053959;
memory[818] = 32'd356728;
memory[819] = 32'd2862806;
memory[820] = 32'd4515797;
memory[821] = 32'd5748720;
memory[822] = 32'd9547084;
memory[823] = 32'd9121308;
memory[824] = 32'd4515334;
memory[825] = 32'd1742698;
memory[826] = 32'd4110991;
memory[827] = 32'd7076376;
memory[828] = 32'd5798898;
memory[829] = 32'd1252715;
memory[830] = 32'd801052;
memory[831] = 32'd2825171;
memory[832] = 32'd5218189;
memory[833] = 32'd5771559;
memory[834] = 32'd752506;
memory[835] = 32'd5554010;
memory[836] = 32'd9709016;
memory[837] = 32'd2178224;
memory[838] = 32'd2173109;
memory[839] = 32'd5816539;
memory[840] = 32'd7490000;
memory[841] = 32'd4333378;
memory[842] = 32'd2058109;
memory[843] = 32'd3945053;
memory[844] = 32'd1955081;
memory[845] = 32'd1489114;
memory[846] = 32'd1671338;
memory[847] = 32'd5405989;
memory[848] = 32'd1059426;
memory[849] = 32'd2028067;
memory[850] = 32'd785147;
memory[851] = 32'd5575223;
memory[852] = 32'd7776787;
memory[853] = 32'd332231;
memory[854] = 32'd4696532;
memory[855] = 32'd2292122;
memory[856] = 32'd4591281;
memory[857] = 32'd1323875;
memory[858] = 32'd1884850;
memory[859] = 32'd390179;
memory[860] = 32'd2576590;
memory[861] = 32'd5202254;
memory[862] = 32'd3215350;
memory[863] = 32'd311131;
memory[864] = 32'd973813;
memory[865] = 32'd3967857;
memory[866] = 32'd8381494;
memory[867] = 32'd3199181;
memory[868] = 32'd6146081;
memory[869] = 32'd554603;
memory[870] = 32'd9015720;
memory[871] = 32'd6152433;
memory[872] = 32'd4887982;
memory[873] = 32'd3590181;
memory[874] = 32'd97487;
memory[875] = 32'd9359415;
memory[876] = 32'd5079296;
memory[877] = 32'd1768825;
memory[878] = 32'd4765404;
memory[879] = 32'd6138722;
memory[880] = 32'd3796892;
memory[881] = 32'd5550551;
memory[882] = 32'd4230297;
memory[883] = 32'd4090032;
memory[884] = 32'd8399134;
memory[885] = 32'd1443181;
memory[886] = 32'd8898506;
memory[887] = 32'd2990415;
memory[888] = 32'd2767057;
memory[889] = 32'd3299708;
memory[890] = 32'd3380595;
memory[891] = 32'd7859999;
memory[892] = 32'd8501962;
memory[893] = 32'd9112297;
memory[894] = 32'd687483;
memory[895] = 32'd9475776;
memory[896] = 32'd3080154;
memory[897] = 32'd9068977;
memory[898] = 32'd5191309;
memory[899] = 32'd1742587;
memory[900] = 32'd2139932;
memory[901] = 32'd6723382;
memory[902] = 32'd7895021;
memory[903] = 32'd9544266;
memory[904] = 32'd313563;
memory[905] = 32'd508860;
memory[906] = 32'd8903682;
memory[907] = 32'd7909211;
memory[908] = 32'd2277685;
memory[909] = 32'd3669086;
memory[910] = 32'd6564285;
memory[911] = 32'd8590930;
memory[912] = 32'd1735990;
memory[913] = 32'd794583;
memory[914] = 32'd5197314;
memory[915] = 32'd2651476;
memory[916] = 32'd4754116;
memory[917] = 32'd4095820;
memory[918] = 32'd5641892;
memory[919] = 32'd37525;
memory[920] = 32'd7395528;
memory[921] = 32'd1538839;
memory[922] = 32'd7897525;
memory[923] = 32'd5897490;
memory[924] = 32'd651136;
memory[925] = 32'd1101360;
memory[926] = 32'd7889618;
memory[927] = 32'd6247643;
memory[928] = 32'd170337;
memory[929] = 32'd3080928;
memory[930] = 32'd506582;
memory[931] = 32'd4826621;
memory[932] = 32'd9804310;
memory[933] = 32'd917955;
memory[934] = 32'd4370888;
memory[935] = 32'd2634225;
memory[936] = 32'd1426815;
memory[937] = 32'd3274570;
memory[938] = 32'd543437;
memory[939] = 32'd6220853;
memory[940] = 32'd9460008;
memory[941] = 32'd7107722;
memory[942] = 32'd4811783;
memory[943] = 32'd3712350;
memory[944] = 32'd418657;
memory[945] = 32'd9097;
memory[946] = 32'd6363827;
memory[947] = 32'd7689126;
memory[948] = 32'd6621269;
memory[949] = 32'd4522071;
memory[950] = 32'd7726651;
memory[951] = 32'd6533149;
memory[952] = 32'd6060910;
memory[953] = 32'd8140528;
memory[954] = 32'd2430639;
memory[955] = 32'd9228398;
memory[956] = 32'd9241888;
memory[957] = 32'd2836610;
memory[958] = 32'd7992393;
memory[959] = 32'd1928577;
memory[960] = 32'd8433890;
memory[961] = 32'd8498976;
memory[962] = 32'd6755199;
memory[963] = 32'd754552;
memory[964] = 32'd9416931;
memory[965] = 32'd1126087;
memory[966] = 32'd3388777;
memory[967] = 32'd3360099;
memory[968] = 32'd4400657;
memory[969] = 32'd6448566;
memory[970] = 32'd9580952;
memory[971] = 32'd6377017;
memory[972] = 32'd6072641;
memory[973] = 32'd4392735;
memory[974] = 32'd89368;
memory[975] = 32'd6491298;
memory[976] = 32'd6918184;
memory[977] = 32'd6453195;
memory[978] = 32'd6696776;
memory[979] = 32'd6055805;
memory[980] = 32'd975266;
memory[981] = 32'd4423428;
memory[982] = 32'd2588954;
memory[983] = 32'd9552528;
memory[984] = 32'd5080308;
memory[985] = 32'd5019593;
memory[986] = 32'd1297278;
memory[987] = 32'd4322197;
memory[988] = 32'd372555;
memory[989] = 32'd9289672;
memory[990] = 32'd6250774;
memory[991] = 32'd8806445;
memory[992] = 32'd305000;
memory[993] = 32'd5522325;
memory[994] = 32'd9560997;
memory[995] = 32'd2238283;
memory[996] = 32'd6648412;
memory[997] = 32'd5466127;
memory[998] = 32'd5598382;
memory[999] = 32'd3565421;
memory[1000] = 32'd1914693;
memory[1001] = 32'd5179334;
memory[1002] = 32'd9942439;
memory[1003] = 32'd7987334;
memory[1004] = 32'd2088421;
memory[1005] = 32'd2548159;
memory[1006] = 32'd6994985;
memory[1007] = 32'd1522957;
memory[1008] = 32'd9001354;
memory[1009] = 32'd3691761;
memory[1010] = 32'd7578762;
memory[1011] = 32'd2492972;
memory[1012] = 32'd631541;
memory[1013] = 32'd167716;
memory[1014] = 32'd4561852;
memory[1015] = 32'd5711850;
memory[1016] = 32'd7703662;
memory[1017] = 32'd8375482;
memory[1018] = 32'd2550399;
memory[1019] = 32'd8076217;
memory[1020] = 32'd7665154;
memory[1021] = 32'd8801173;
memory[1022] = 32'd9399015;
memory[1023] = 32'd486506;
memory[1024] = 32'd6839851;
memory[1025] = 32'd1476364;
memory[1026] = 32'd2724790;
memory[1027] = 32'd3488263;
memory[1028] = 32'd6942491;
memory[1029] = 32'd8323172;
memory[1030] = 32'd9570037;
memory[1031] = 32'd1373537;
memory[1032] = 32'd6018859;
memory[1033] = 32'd2028828;
memory[1034] = 32'd9360871;
memory[1035] = 32'd8107280;
memory[1036] = 32'd4576987;
memory[1037] = 32'd6355856;
memory[1038] = 32'd2146590;
memory[1039] = 32'd3578341;
memory[1040] = 32'd2563970;
memory[1041] = 32'd9725352;
memory[1042] = 32'd8587665;
memory[1043] = 32'd3195511;
memory[1044] = 32'd9893069;
memory[1045] = 32'd3149517;
memory[1046] = 32'd8907361;
memory[1047] = 32'd113083;
memory[1048] = 32'd4041351;
memory[1049] = 32'd3974112;
memory[1050] = 32'd8189300;
memory[1051] = 32'd1706506;
memory[1052] = 32'd5291638;
memory[1053] = 32'd104667;
memory[1054] = 32'd4709364;
memory[1055] = 32'd2131489;
memory[1056] = 32'd1581032;
memory[1057] = 32'd7434154;
memory[1058] = 32'd8136104;
memory[1059] = 32'd1039875;
memory[1060] = 32'd8273679;
memory[1061] = 32'd7706141;
memory[1062] = 32'd2413412;
memory[1063] = 32'd4292538;
memory[1064] = 32'd9734969;
memory[1065] = 32'd4290636;
memory[1066] = 32'd4916170;
memory[1067] = 32'd4311956;
memory[1068] = 32'd3162844;
memory[1069] = 32'd7062760;
memory[1070] = 32'd406649;
memory[1071] = 32'd5726814;
memory[1072] = 32'd9304465;
memory[1073] = 32'd8994314;
memory[1074] = 32'd8922326;
memory[1075] = 32'd1713886;
memory[1076] = 32'd4660183;
memory[1077] = 32'd346039;
memory[1078] = 32'd1826969;
memory[1079] = 32'd8701535;
memory[1080] = 32'd4320152;
memory[1081] = 32'd2532621;
memory[1082] = 32'd2924393;
memory[1083] = 32'd9611790;
memory[1084] = 32'd2637289;
memory[1085] = 32'd150109;
memory[1086] = 32'd4259631;
memory[1087] = 32'd6734673;
memory[1088] = 32'd7584264;
memory[1089] = 32'd2395735;
memory[1090] = 32'd7774548;
memory[1091] = 32'd8374295;
memory[1092] = 32'd101877;
memory[1093] = 32'd2704313;
memory[1094] = 32'd2666833;
memory[1095] = 32'd2353198;
memory[1096] = 32'd6994949;
memory[1097] = 32'd99355;
memory[1098] = 32'd6665155;
memory[1099] = 32'd157793;
memory[1100] = 32'd9678468;
memory[1101] = 32'd9588156;
memory[1102] = 32'd8400960;
memory[1103] = 32'd8982933;
memory[1104] = 32'd1098823;
memory[1105] = 32'd7323286;
memory[1106] = 32'd3213171;
memory[1107] = 32'd8275358;
memory[1108] = 32'd185677;
memory[1109] = 32'd5040140;
memory[1110] = 32'd9493245;
memory[1111] = 32'd7022181;
memory[1112] = 32'd7572761;
memory[1113] = 32'd4933990;
memory[1114] = 32'd9150323;
memory[1115] = 32'd210050;
memory[1116] = 32'd5084100;
memory[1117] = 32'd3409954;
memory[1118] = 32'd9461075;
memory[1119] = 32'd2668364;
memory[1120] = 32'd8322042;
memory[1121] = 32'd7235624;
memory[1122] = 32'd1042659;
memory[1123] = 32'd8423919;
memory[1124] = 32'd2456289;
memory[1125] = 32'd6225844;
memory[1126] = 32'd3293469;
memory[1127] = 32'd9451238;
memory[1128] = 32'd8841551;
memory[1129] = 32'd2474976;
memory[1130] = 32'd2125383;
memory[1131] = 32'd8520019;
memory[1132] = 32'd2063133;
memory[1133] = 32'd526343;
memory[1134] = 32'd19304;
memory[1135] = 32'd3161956;
memory[1136] = 32'd365981;
memory[1137] = 32'd3232475;
memory[1138] = 32'd3953666;
memory[1139] = 32'd3068011;
memory[1140] = 32'd788967;
memory[1141] = 32'd3446912;
memory[1142] = 32'd90192;
memory[1143] = 32'd8361729;
memory[1144] = 32'd8380902;
memory[1145] = 32'd1756868;
memory[1146] = 32'd1088131;
memory[1147] = 32'd3465002;
memory[1148] = 32'd7683174;
memory[1149] = 32'd549207;
memory[1150] = 32'd8649718;
memory[1151] = 32'd6005216;
memory[1152] = 32'd301183;
memory[1153] = 32'd9692377;
memory[1154] = 32'd6945487;
memory[1155] = 32'd2757472;
memory[1156] = 32'd8434573;
memory[1157] = 32'd238957;
memory[1158] = 32'd4725062;
memory[1159] = 32'd7276125;
memory[1160] = 32'd2713933;
memory[1161] = 32'd9366797;
memory[1162] = 32'd8312496;
memory[1163] = 32'd7293418;
memory[1164] = 32'd9893141;
memory[1165] = 32'd848153;
memory[1166] = 32'd2971726;
memory[1167] = 32'd2775474;
memory[1168] = 32'd6596980;
memory[1169] = 32'd6925393;
memory[1170] = 32'd5843485;
memory[1171] = 32'd7385948;
memory[1172] = 32'd372305;
memory[1173] = 32'd8450030;
memory[1174] = 32'd8264029;
memory[1175] = 32'd1269559;
memory[1176] = 32'd206898;
memory[1177] = 32'd9352160;
memory[1178] = 32'd4734562;
memory[1179] = 32'd406424;
memory[1180] = 32'd2417719;
memory[1181] = 32'd3384280;
memory[1182] = 32'd6411641;
memory[1183] = 32'd2718902;
memory[1184] = 32'd5593010;
memory[1185] = 32'd5873480;
memory[1186] = 32'd7992726;
memory[1187] = 32'd4027583;
memory[1188] = 32'd8628789;
memory[1189] = 32'd5234140;
memory[1190] = 32'd1303708;
memory[1191] = 32'd1342723;
memory[1192] = 32'd4600938;
memory[1193] = 32'd2132557;
memory[1194] = 32'd1152493;
memory[1195] = 32'd7010431;
memory[1196] = 32'd2980710;
memory[1197] = 32'd4124220;
memory[1198] = 32'd9785905;
memory[1199] = 32'd9577690;
memory[1200] = 32'd1049613;
memory[1201] = 32'd5629391;
memory[1202] = 32'd6963638;
memory[1203] = 32'd3938270;
memory[1204] = 32'd4079421;
memory[1205] = 32'd5227667;
memory[1206] = 32'd5207829;
memory[1207] = 32'd6802671;
memory[1208] = 32'd7096180;
memory[1209] = 32'd2458743;
memory[1210] = 32'd7209095;
memory[1211] = 32'd9513899;
memory[1212] = 32'd5843024;
memory[1213] = 32'd6137088;
memory[1214] = 32'd4749154;
memory[1215] = 32'd3952386;
memory[1216] = 32'd2010569;
memory[1217] = 32'd5258232;
memory[1218] = 32'd7979969;
memory[1219] = 32'd3155710;
memory[1220] = 32'd492373;
memory[1221] = 32'd1800030;
memory[1222] = 32'd4498433;
memory[1223] = 32'd7609663;
memory[1224] = 32'd3932587;
memory[1225] = 32'd8167279;
memory[1226] = 32'd4620094;
memory[1227] = 32'd9429649;
memory[1228] = 32'd2291499;
memory[1229] = 32'd6922351;
memory[1230] = 32'd9007339;
memory[1231] = 32'd5857464;
memory[1232] = 32'd2551742;
memory[1233] = 32'd8487330;
memory[1234] = 32'd2312086;
memory[1235] = 32'd9147515;
memory[1236] = 32'd6231349;
memory[1237] = 32'd7519915;
memory[1238] = 32'd5950186;
memory[1239] = 32'd5843881;
memory[1240] = 32'd2495011;
memory[1241] = 32'd5675634;
memory[1242] = 32'd7874133;
memory[1243] = 32'd854387;
memory[1244] = 32'd1812722;
memory[1245] = 32'd2623287;
memory[1246] = 32'd4806773;
memory[1247] = 32'd6339643;
memory[1248] = 32'd7881519;
memory[1249] = 32'd2786742;
memory[1250] = 32'd9495354;
memory[1251] = 32'd890244;
memory[1252] = 32'd7103124;
memory[1253] = 32'd6510139;
memory[1254] = 32'd1016259;
memory[1255] = 32'd3552063;
memory[1256] = 32'd4677418;
memory[1257] = 32'd5636353;
memory[1258] = 32'd2981712;
memory[1259] = 32'd9485269;
memory[1260] = 32'd2558705;
memory[1261] = 32'd4505404;
memory[1262] = 32'd5342733;
memory[1263] = 32'd7626799;
memory[1264] = 32'd2992734;
memory[1265] = 32'd7654819;
memory[1266] = 32'd6774315;
memory[1267] = 32'd1740435;
memory[1268] = 32'd7691087;
memory[1269] = 32'd5240853;
memory[1270] = 32'd100669;
memory[1271] = 32'd2702450;
memory[1272] = 32'd916487;
memory[1273] = 32'd7974802;
memory[1274] = 32'd3556837;
memory[1275] = 32'd5245562;
memory[1276] = 32'd598089;
memory[1277] = 32'd8363610;
memory[1278] = 32'd1585205;
memory[1279] = 32'd995960;
memory[1280] = 32'd3666704;
memory[1281] = 32'd3596911;
memory[1282] = 32'd4402557;
memory[1283] = 32'd769829;
memory[1284] = 32'd2623403;
memory[1285] = 32'd5418816;
memory[1286] = 32'd4321892;
memory[1287] = 32'd7300821;
memory[1288] = 32'd3571522;
memory[1289] = 32'd7303605;
memory[1290] = 32'd9302443;
memory[1291] = 32'd8646579;
memory[1292] = 32'd4325361;
memory[1293] = 32'd7161528;
memory[1294] = 32'd6273378;
memory[1295] = 32'd9834447;
memory[1296] = 32'd7332700;
memory[1297] = 32'd5564045;
memory[1298] = 32'd1574882;
memory[1299] = 32'd5023787;
memory[1300] = 32'd804899;
memory[1301] = 32'd1675551;
memory[1302] = 32'd242589;
memory[1303] = 32'd1721386;
memory[1304] = 32'd9650353;
memory[1305] = 32'd3799426;
memory[1306] = 32'd6966948;
memory[1307] = 32'd2764794;
memory[1308] = 32'd2163036;
memory[1309] = 32'd1068506;
memory[1310] = 32'd6277107;
memory[1311] = 32'd8346092;
memory[1312] = 32'd4665417;
memory[1313] = 32'd679664;
memory[1314] = 32'd9115921;
memory[1315] = 32'd7288820;
memory[1316] = 32'd6098480;
memory[1317] = 32'd5954166;
memory[1318] = 32'd7105994;
memory[1319] = 32'd2186354;
memory[1320] = 32'd5774123;
memory[1321] = 32'd6408437;
memory[1322] = 32'd832933;
memory[1323] = 32'd99484;
memory[1324] = 32'd6086317;
memory[1325] = 32'd7106312;
memory[1326] = 32'd9933931;
memory[1327] = 32'd3419017;
memory[1328] = 32'd5186709;
memory[1329] = 32'd4025165;
memory[1330] = 32'd959156;
memory[1331] = 32'd5991608;
memory[1332] = 32'd8217069;
memory[1333] = 32'd1201745;
memory[1334] = 32'd7712995;
memory[1335] = 32'd7867422;
memory[1336] = 32'd5001171;
memory[1337] = 32'd7196295;
memory[1338] = 32'd3148569;
memory[1339] = 32'd9680559;
memory[1340] = 32'd8264801;
memory[1341] = 32'd9425676;
memory[1342] = 32'd8026652;
memory[1343] = 32'd5446571;
memory[1344] = 32'd105340;
memory[1345] = 32'd9658925;
memory[1346] = 32'd5251743;
memory[1347] = 32'd8720172;
memory[1348] = 32'd5613091;
memory[1349] = 32'd4874089;
memory[1350] = 32'd906527;
memory[1351] = 32'd3903566;
memory[1352] = 32'd3798878;
memory[1353] = 32'd4255812;
memory[1354] = 32'd4003050;
memory[1355] = 32'd9885196;
memory[1356] = 32'd1362124;
memory[1357] = 32'd6453333;
memory[1358] = 32'd3304213;
memory[1359] = 32'd9065186;
memory[1360] = 32'd478499;
memory[1361] = 32'd4263370;
memory[1362] = 32'd5056794;
memory[1363] = 32'd8695568;
memory[1364] = 32'd5465115;
memory[1365] = 32'd5286141;
memory[1366] = 32'd9079342;
memory[1367] = 32'd2982639;
memory[1368] = 32'd2482437;
memory[1369] = 32'd4744263;
memory[1370] = 32'd2663198;
memory[1371] = 32'd3263590;
memory[1372] = 32'd4169939;
memory[1373] = 32'd3206202;
memory[1374] = 32'd1226513;
memory[1375] = 32'd6791631;
memory[1376] = 32'd2865128;
memory[1377] = 32'd6478257;
memory[1378] = 32'd5511804;
memory[1379] = 32'd994571;
memory[1380] = 32'd1352346;
memory[1381] = 32'd8934683;
memory[1382] = 32'd4898138;
memory[1383] = 32'd5151225;
memory[1384] = 32'd3190495;
memory[1385] = 32'd1417540;
memory[1386] = 32'd5036421;
memory[1387] = 32'd7068972;
memory[1388] = 32'd387226;
memory[1389] = 32'd8340634;
memory[1390] = 32'd6134158;
memory[1391] = 32'd865725;
memory[1392] = 32'd5120356;
memory[1393] = 32'd1190952;
memory[1394] = 32'd2077645;
memory[1395] = 32'd585472;
memory[1396] = 32'd8993446;
memory[1397] = 32'd3673339;
memory[1398] = 32'd3568111;
memory[1399] = 32'd1475883;
memory[1400] = 32'd8417603;
memory[1401] = 32'd8747661;
memory[1402] = 32'd7255825;
memory[1403] = 32'd2587542;
memory[1404] = 32'd4470216;
memory[1405] = 32'd8482339;
memory[1406] = 32'd9379174;
memory[1407] = 32'd7335344;
memory[1408] = 32'd4960596;
memory[1409] = 32'd7407330;
memory[1410] = 32'd846267;
memory[1411] = 32'd8829294;
memory[1412] = 32'd6342013;
memory[1413] = 32'd8260757;
memory[1414] = 32'd3980519;
memory[1415] = 32'd2048860;
memory[1416] = 32'd2194650;
memory[1417] = 32'd1533292;
memory[1418] = 32'd9117832;
memory[1419] = 32'd2581876;
memory[1420] = 32'd2390279;
memory[1421] = 32'd5251990;
memory[1422] = 32'd5963953;
memory[1423] = 32'd7510635;
memory[1424] = 32'd8959295;
memory[1425] = 32'd8041598;
memory[1426] = 32'd8096107;
memory[1427] = 32'd7952741;
memory[1428] = 32'd1714937;
memory[1429] = 32'd4180570;
memory[1430] = 32'd1944976;
memory[1431] = 32'd132540;
memory[1432] = 32'd5444584;
memory[1433] = 32'd9200801;
memory[1434] = 32'd2720083;
memory[1435] = 32'd9914800;
memory[1436] = 32'd199492;
memory[1437] = 32'd4615609;
memory[1438] = 32'd9766496;
memory[1439] = 32'd7676440;
memory[1440] = 32'd2022939;
memory[1441] = 32'd612763;
memory[1442] = 32'd6505735;
memory[1443] = 32'd881304;
memory[1444] = 32'd1389873;
memory[1445] = 32'd3002606;
memory[1446] = 32'd2930164;
memory[1447] = 32'd3584523;
memory[1448] = 32'd7052251;
memory[1449] = 32'd4564349;
memory[1450] = 32'd8682751;
memory[1451] = 32'd9442530;
memory[1452] = 32'd9816339;
memory[1453] = 32'd4646704;
memory[1454] = 32'd6953165;
memory[1455] = 32'd1291986;
memory[1456] = 32'd2688302;
memory[1457] = 32'd7565625;
memory[1458] = 32'd1761079;
memory[1459] = 32'd6919591;
memory[1460] = 32'd4262547;
memory[1461] = 32'd6222407;
memory[1462] = 32'd9568484;
memory[1463] = 32'd9707131;
memory[1464] = 32'd7939561;
memory[1465] = 32'd4804919;
memory[1466] = 32'd9621931;
memory[1467] = 32'd8139053;
memory[1468] = 32'd9420528;
memory[1469] = 32'd9388427;
memory[1470] = 32'd5815494;
memory[1471] = 32'd3959819;
memory[1472] = 32'd2517543;
memory[1473] = 32'd4837581;
memory[1474] = 32'd4841123;
memory[1475] = 32'd6423768;
memory[1476] = 32'd7840187;
memory[1477] = 32'd287639;
memory[1478] = 32'd2524643;
memory[1479] = 32'd4892438;
memory[1480] = 32'd4851988;
memory[1481] = 32'd1207394;
memory[1482] = 32'd6851320;
memory[1483] = 32'd7184680;
memory[1484] = 32'd5854098;
memory[1485] = 32'd3804486;
memory[1486] = 32'd993018;
memory[1487] = 32'd1058752;
memory[1488] = 32'd3886463;
memory[1489] = 32'd2754098;
memory[1490] = 32'd494695;
memory[1491] = 32'd8149010;
memory[1492] = 32'd8976505;
memory[1493] = 32'd63179;
memory[1494] = 32'd7856142;
memory[1495] = 32'd6916066;
memory[1496] = 32'd4868098;
memory[1497] = 32'd9994425;
memory[1498] = 32'd7571472;
memory[1499] = 32'd6804978;
memory[1500] = 32'd9382853;
memory[1501] = 32'd3386966;
memory[1502] = 32'd764797;
memory[1503] = 32'd4416748;
memory[1504] = 32'd8224547;
memory[1505] = 32'd8122272;
memory[1506] = 32'd840516;
memory[1507] = 32'd8581086;
memory[1508] = 32'd8409912;
memory[1509] = 32'd3365159;
memory[1510] = 32'd5989877;
memory[1511] = 32'd3261900;
memory[1512] = 32'd4572553;
memory[1513] = 32'd2841197;
memory[1514] = 32'd2962932;
memory[1515] = 32'd2943003;
memory[1516] = 32'd9162035;
memory[1517] = 32'd3955951;
memory[1518] = 32'd6518107;
memory[1519] = 32'd3048498;
memory[1520] = 32'd6710049;
memory[1521] = 32'd9529154;
memory[1522] = 32'd3713861;
memory[1523] = 32'd8202906;
memory[1524] = 32'd9592334;
memory[1525] = 32'd1570003;
memory[1526] = 32'd7635325;
memory[1527] = 32'd6976784;
memory[1528] = 32'd1564428;
memory[1529] = 32'd5206797;
memory[1530] = 32'd3781763;
memory[1531] = 32'd3463633;
memory[1532] = 32'd1110115;
memory[1533] = 32'd4546560;
memory[1534] = 32'd7880381;
memory[1535] = 32'd1851014;
memory[1536] = 32'd5185185;
memory[1537] = 32'd8720897;
memory[1538] = 32'd432100;
memory[1539] = 32'd3595097;
memory[1540] = 32'd4602408;
memory[1541] = 32'd8938329;
memory[1542] = 32'd9373349;
memory[1543] = 32'd1691313;
memory[1544] = 32'd4295879;
memory[1545] = 32'd4852634;
memory[1546] = 32'd4634316;
memory[1547] = 32'd3457914;
memory[1548] = 32'd8808585;
memory[1549] = 32'd3668775;
memory[1550] = 32'd9022765;
memory[1551] = 32'd8034986;
memory[1552] = 32'd3197930;
memory[1553] = 32'd2736626;
memory[1554] = 32'd6237892;
memory[1555] = 32'd5306616;
memory[1556] = 32'd4306629;
memory[1557] = 32'd6389569;
memory[1558] = 32'd4799752;
memory[1559] = 32'd8387409;
memory[1560] = 32'd1596366;
memory[1561] = 32'd8581515;
memory[1562] = 32'd4367395;
memory[1563] = 32'd5222833;
memory[1564] = 32'd5644428;
memory[1565] = 32'd2247776;
memory[1566] = 32'd7073847;
memory[1567] = 32'd829613;
memory[1568] = 32'd3485026;
memory[1569] = 32'd22300;
memory[1570] = 32'd6941062;
memory[1571] = 32'd603786;
memory[1572] = 32'd8960629;
memory[1573] = 32'd8830763;
memory[1574] = 32'd2295100;
memory[1575] = 32'd3256508;
memory[1576] = 32'd3683397;
memory[1577] = 32'd6929416;
memory[1578] = 32'd9230775;
memory[1579] = 32'd2491982;
memory[1580] = 32'd3114544;
memory[1581] = 32'd8253540;
memory[1582] = 32'd3043320;
memory[1583] = 32'd8828826;
memory[1584] = 32'd3506518;
memory[1585] = 32'd1797565;
memory[1586] = 32'd6651794;
memory[1587] = 32'd329499;
memory[1588] = 32'd8187134;
memory[1589] = 32'd1451546;
memory[1590] = 32'd8716908;
memory[1591] = 32'd2299853;
memory[1592] = 32'd33062;
memory[1593] = 32'd3084303;
memory[1594] = 32'd7522686;
memory[1595] = 32'd8193842;
memory[1596] = 32'd7848432;
memory[1597] = 32'd4596534;
memory[1598] = 32'd1539807;
memory[1599] = 32'd3849810;
memory[1600] = 32'd4618834;
memory[1601] = 32'd8480869;
memory[1602] = 32'd4453596;
memory[1603] = 32'd6095815;
memory[1604] = 32'd9827984;
memory[1605] = 32'd6748696;
memory[1606] = 32'd9352324;
memory[1607] = 32'd3511382;
memory[1608] = 32'd6194465;
memory[1609] = 32'd1099451;
memory[1610] = 32'd8519716;
memory[1611] = 32'd1825361;
memory[1612] = 32'd1869343;
memory[1613] = 32'd1563037;
memory[1614] = 32'd654187;
memory[1615] = 32'd5375861;
memory[1616] = 32'd3360602;
memory[1617] = 32'd7305981;
memory[1618] = 32'd5705360;
memory[1619] = 32'd4064088;
memory[1620] = 32'd1273879;
memory[1621] = 32'd6938620;
memory[1622] = 32'd6363941;
memory[1623] = 32'd3823293;
memory[1624] = 32'd22924;
memory[1625] = 32'd3886628;
memory[1626] = 32'd2017135;
memory[1627] = 32'd387708;
memory[1628] = 32'd8483162;
memory[1629] = 32'd3556942;
memory[1630] = 32'd6753870;
memory[1631] = 32'd3101996;
memory[1632] = 32'd4554163;
memory[1633] = 32'd1207466;
memory[1634] = 32'd9197811;
memory[1635] = 32'd6898500;
memory[1636] = 32'd472515;
memory[1637] = 32'd1066487;
memory[1638] = 32'd2926234;
memory[1639] = 32'd9183332;
memory[1640] = 32'd4682290;
memory[1641] = 32'd1445950;
memory[1642] = 32'd1008693;
memory[1643] = 32'd6551633;
memory[1644] = 32'd5525339;
memory[1645] = 32'd1662880;
memory[1646] = 32'd1927494;
memory[1647] = 32'd1402293;
memory[1648] = 32'd1485213;
memory[1649] = 32'd7632854;
memory[1650] = 32'd5466382;
memory[1651] = 32'd5275444;
memory[1652] = 32'd4571475;
memory[1653] = 32'd1830323;
memory[1654] = 32'd9098738;
memory[1655] = 32'd7110751;
memory[1656] = 32'd5716951;
memory[1657] = 32'd1115873;
memory[1658] = 32'd14811;
memory[1659] = 32'd6716465;
memory[1660] = 32'd7189168;
memory[1661] = 32'd6768681;
memory[1662] = 32'd2334813;
memory[1663] = 32'd4259683;
memory[1664] = 32'd492499;
memory[1665] = 32'd4048977;
memory[1666] = 32'd3674535;
memory[1667] = 32'd965014;
memory[1668] = 32'd5115464;
memory[1669] = 32'd6600769;
memory[1670] = 32'd148346;
memory[1671] = 32'd2314107;
memory[1672] = 32'd563072;
memory[1673] = 32'd3673391;
memory[1674] = 32'd8865740;
memory[1675] = 32'd6088411;
memory[1676] = 32'd7852623;
memory[1677] = 32'd3309587;
memory[1678] = 32'd7057;
memory[1679] = 32'd9337836;
memory[1680] = 32'd3458793;
memory[1681] = 32'd5473439;
memory[1682] = 32'd4613281;
memory[1683] = 32'd546620;
memory[1684] = 32'd9820114;
memory[1685] = 32'd6228371;
memory[1686] = 32'd7657371;
memory[1687] = 32'd8053418;
memory[1688] = 32'd9860596;
memory[1689] = 32'd188534;
memory[1690] = 32'd4769883;
memory[1691] = 32'd7049764;
memory[1692] = 32'd9473567;
memory[1693] = 32'd7104697;
memory[1694] = 32'd3825800;
memory[1695] = 32'd9966067;
memory[1696] = 32'd1153674;
memory[1697] = 32'd7500335;
memory[1698] = 32'd3447433;
memory[1699] = 32'd8785490;
memory[1700] = 32'd6617457;
memory[1701] = 32'd6112132;
memory[1702] = 32'd3615949;
memory[1703] = 32'd7180529;
memory[1704] = 32'd9785523;
memory[1705] = 32'd2481690;
memory[1706] = 32'd5785292;
memory[1707] = 32'd7638147;
memory[1708] = 32'd8307629;
memory[1709] = 32'd5792349;
memory[1710] = 32'd9492335;
memory[1711] = 32'd1766422;
memory[1712] = 32'd3782140;
memory[1713] = 32'd6621968;
memory[1714] = 32'd2313043;
memory[1715] = 32'd3602255;
memory[1716] = 32'd2850339;
memory[1717] = 32'd2486766;
memory[1718] = 32'd4172025;
memory[1719] = 32'd2710936;
memory[1720] = 32'd5191653;
memory[1721] = 32'd1458260;
memory[1722] = 32'd2277052;
memory[1723] = 32'd4665220;
memory[1724] = 32'd8562957;
memory[1725] = 32'd8619204;
memory[1726] = 32'd4631287;
memory[1727] = 32'd2232983;
memory[1728] = 32'd6119540;
memory[1729] = 32'd8078721;
memory[1730] = 32'd3534826;
memory[1731] = 32'd2736997;
memory[1732] = 32'd6707205;
memory[1733] = 32'd9667127;
memory[1734] = 32'd2433878;
memory[1735] = 32'd6492728;
memory[1736] = 32'd4665169;
memory[1737] = 32'd8219170;
memory[1738] = 32'd6647227;
memory[1739] = 32'd2972798;
memory[1740] = 32'd4011520;
memory[1741] = 32'd6139563;
memory[1742] = 32'd4739221;
memory[1743] = 32'd7793660;
memory[1744] = 32'd5277883;
memory[1745] = 32'd9568616;
memory[1746] = 32'd3912267;
memory[1747] = 32'd8128223;
memory[1748] = 32'd2055382;
memory[1749] = 32'd8084292;
memory[1750] = 32'd3355511;
memory[1751] = 32'd7247035;
memory[1752] = 32'd9542553;
memory[1753] = 32'd5632563;
memory[1754] = 32'd4428608;
memory[1755] = 32'd621862;
memory[1756] = 32'd4251768;
memory[1757] = 32'd9059895;
memory[1758] = 32'd5371198;
memory[1759] = 32'd2887660;
memory[1760] = 32'd9654968;
memory[1761] = 32'd1422376;
memory[1762] = 32'd8141009;
memory[1763] = 32'd6362173;
memory[1764] = 32'd1089503;
memory[1765] = 32'd574887;
memory[1766] = 32'd5371254;
memory[1767] = 32'd5754673;
memory[1768] = 32'd8794057;
memory[1769] = 32'd2018481;
memory[1770] = 32'd1243823;
memory[1771] = 32'd5321929;
memory[1772] = 32'd674396;
memory[1773] = 32'd5983044;
memory[1774] = 32'd5631942;
memory[1775] = 32'd5952280;
memory[1776] = 32'd8068012;
memory[1777] = 32'd9544209;
memory[1778] = 32'd6596855;
memory[1779] = 32'd2639747;
memory[1780] = 32'd144854;
memory[1781] = 32'd9952366;
memory[1782] = 32'd2403134;
memory[1783] = 32'd2203759;
memory[1784] = 32'd8101281;
memory[1785] = 32'd6831742;
memory[1786] = 32'd5341973;
memory[1787] = 32'd4869401;
memory[1788] = 32'd5891638;
memory[1789] = 32'd713171;
memory[1790] = 32'd273413;
memory[1791] = 32'd8062958;
memory[1792] = 32'd4651899;
memory[1793] = 32'd8414422;
memory[1794] = 32'd6941484;
memory[1795] = 32'd8257755;
memory[1796] = 32'd1505661;
memory[1797] = 32'd4829090;
memory[1798] = 32'd6528780;
memory[1799] = 32'd2816071;
memory[1800] = 32'd9363923;
memory[1801] = 32'd7772603;
memory[1802] = 32'd8138000;
memory[1803] = 32'd38320;
memory[1804] = 32'd6272000;
memory[1805] = 32'd3769942;
memory[1806] = 32'd8506952;
memory[1807] = 32'd4340012;
memory[1808] = 32'd5830504;
memory[1809] = 32'd5103807;
memory[1810] = 32'd6979759;
memory[1811] = 32'd5975358;
memory[1812] = 32'd7572525;
memory[1813] = 32'd9382894;
memory[1814] = 32'd8179117;
memory[1815] = 32'd8190158;
memory[1816] = 32'd6214636;
memory[1817] = 32'd3521090;
memory[1818] = 32'd3059560;
memory[1819] = 32'd4622626;
memory[1820] = 32'd6750614;
memory[1821] = 32'd3332973;
memory[1822] = 32'd5201937;
memory[1823] = 32'd3918865;
memory[1824] = 32'd4263748;
memory[1825] = 32'd2143421;
memory[1826] = 32'd2176620;
memory[1827] = 32'd5769409;
memory[1828] = 32'd9488863;
memory[1829] = 32'd8705400;
memory[1830] = 32'd1101832;
memory[1831] = 32'd8852786;
memory[1832] = 32'd6478004;
memory[1833] = 32'd9239833;
memory[1834] = 32'd1407458;
memory[1835] = 32'd5266356;
memory[1836] = 32'd5526127;
memory[1837] = 32'd9914410;
memory[1838] = 32'd9606368;
memory[1839] = 32'd1356631;
memory[1840] = 32'd7534569;
memory[1841] = 32'd6586128;
memory[1842] = 32'd9848341;
memory[1843] = 32'd7623446;
memory[1844] = 32'd8485374;
memory[1845] = 32'd8027458;
memory[1846] = 32'd5813605;
memory[1847] = 32'd4700010;
memory[1848] = 32'd4064901;
memory[1849] = 32'd8873165;
memory[1850] = 32'd1838989;
memory[1851] = 32'd3331867;
memory[1852] = 32'd4722490;
memory[1853] = 32'd7040926;
memory[1854] = 32'd7250732;
memory[1855] = 32'd8986238;
memory[1856] = 32'd1700699;
memory[1857] = 32'd1943705;
memory[1858] = 32'd7272000;
memory[1859] = 32'd1189562;
memory[1860] = 32'd3165457;
memory[1861] = 32'd8373832;
memory[1862] = 32'd42348;
memory[1863] = 32'd9643461;
memory[1864] = 32'd130017;
memory[1865] = 32'd1449807;
memory[1866] = 32'd7426169;
memory[1867] = 32'd8172497;
memory[1868] = 32'd3880569;
memory[1869] = 32'd7032538;
memory[1870] = 32'd9529128;
memory[1871] = 32'd1415139;
memory[1872] = 32'd6135018;
memory[1873] = 32'd9377470;
memory[1874] = 32'd9038585;
memory[1875] = 32'd4620392;
memory[1876] = 32'd9921280;
memory[1877] = 32'd7368542;
memory[1878] = 32'd1836754;
memory[1879] = 32'd6502533;
memory[1880] = 32'd6241707;
memory[1881] = 32'd3675743;
memory[1882] = 32'd9834400;
memory[1883] = 32'd3480550;
memory[1884] = 32'd3233021;
memory[1885] = 32'd9601485;
memory[1886] = 32'd2466788;
memory[1887] = 32'd4933720;
memory[1888] = 32'd1545190;
memory[1889] = 32'd2255140;
memory[1890] = 32'd8639634;
memory[1891] = 32'd4710647;
memory[1892] = 32'd3145325;
memory[1893] = 32'd8681983;
memory[1894] = 32'd6870461;
memory[1895] = 32'd5791694;
memory[1896] = 32'd2648142;
memory[1897] = 32'd4296630;
memory[1898] = 32'd3964191;
memory[1899] = 32'd9045063;
memory[1900] = 32'd3845520;
memory[1901] = 32'd3493320;
memory[1902] = 32'd2976554;
memory[1903] = 32'd9980538;
memory[1904] = 32'd5387142;
memory[1905] = 32'd4531492;
memory[1906] = 32'd4600930;
memory[1907] = 32'd5308422;
memory[1908] = 32'd1900034;
memory[1909] = 32'd6437685;
memory[1910] = 32'd4327308;
memory[1911] = 32'd658094;
memory[1912] = 32'd2629780;
memory[1913] = 32'd4161708;
memory[1914] = 32'd4138644;
memory[1915] = 32'd5862802;
memory[1916] = 32'd6279545;
memory[1917] = 32'd9121784;
memory[1918] = 32'd796522;
memory[1919] = 32'd341087;
memory[1920] = 32'd1376925;
memory[1921] = 32'd9436157;
memory[1922] = 32'd5051735;
memory[1923] = 32'd7038602;
memory[1924] = 32'd634492;
memory[1925] = 32'd4438548;
memory[1926] = 32'd2830296;
memory[1927] = 32'd5798986;
memory[1928] = 32'd1251530;
memory[1929] = 32'd9310840;
memory[1930] = 32'd4844049;
memory[1931] = 32'd5097051;
memory[1932] = 32'd5320512;
memory[1933] = 32'd336956;
memory[1934] = 32'd5077589;
memory[1935] = 32'd707654;
memory[1936] = 32'd4868448;
memory[1937] = 32'd2194872;
memory[1938] = 32'd8532428;
memory[1939] = 32'd6768482;
memory[1940] = 32'd8632557;
memory[1941] = 32'd5376088;
memory[1942] = 32'd7426576;
memory[1943] = 32'd1262337;
memory[1944] = 32'd9537797;
memory[1945] = 32'd1565220;
memory[1946] = 32'd7125139;
memory[1947] = 32'd8333694;
memory[1948] = 32'd687005;
memory[1949] = 32'd438014;
memory[1950] = 32'd8674782;
memory[1951] = 32'd4580282;
memory[1952] = 32'd2390523;
memory[1953] = 32'd6242869;
memory[1954] = 32'd4135236;
memory[1955] = 32'd3025015;
memory[1956] = 32'd681417;
memory[1957] = 32'd9481884;
memory[1958] = 32'd1340353;
memory[1959] = 32'd4449299;
memory[1960] = 32'd8792724;
memory[1961] = 32'd8700754;
memory[1962] = 32'd9546350;
memory[1963] = 32'd4113236;
memory[1964] = 32'd9037710;
memory[1965] = 32'd7140292;
memory[1966] = 32'd7337242;
memory[1967] = 32'd3906158;
memory[1968] = 32'd9335164;
memory[1969] = 32'd8386023;
memory[1970] = 32'd674641;
memory[1971] = 32'd7967721;
memory[1972] = 32'd3762111;
memory[1973] = 32'd617569;
memory[1974] = 32'd1746410;
memory[1975] = 32'd5816260;
memory[1976] = 32'd2182790;
memory[1977] = 32'd1387902;
memory[1978] = 32'd4149955;
memory[1979] = 32'd5386147;
memory[1980] = 32'd1825916;
memory[1981] = 32'd5341089;
memory[1982] = 32'd2482781;
memory[1983] = 32'd4216439;
memory[1984] = 32'd1583958;
memory[1985] = 32'd6618017;
memory[1986] = 32'd9757806;
memory[1987] = 32'd2265375;
memory[1988] = 32'd6099901;
memory[1989] = 32'd3614511;
memory[1990] = 32'd6714674;
memory[1991] = 32'd7408978;
memory[1992] = 32'd2315265;
memory[1993] = 32'd8777377;
memory[1994] = 32'd4038566;
memory[1995] = 32'd1352976;
memory[1996] = 32'd5917669;
memory[1997] = 32'd3892161;
memory[1998] = 32'd5259134;
memory[1999] = 32'd5252833;
memory[2000] = 32'd4794536;
memory[2001] = 32'd8450127;
memory[2002] = 32'd5736906;
memory[2003] = 32'd1072999;
memory[2004] = 32'd9067697;
memory[2005] = 32'd7483316;
memory[2006] = 32'd6889260;
memory[2007] = 32'd3766839;
memory[2008] = 32'd1387570;
memory[2009] = 32'd3555567;
memory[2010] = 32'd9152986;
memory[2011] = 32'd3213486;
memory[2012] = 32'd1413008;
memory[2013] = 32'd1635767;
memory[2014] = 32'd9946277;
memory[2015] = 32'd2996966;
memory[2016] = 32'd770136;
memory[2017] = 32'd2220435;
memory[2018] = 32'd7778693;
memory[2019] = 32'd6870037;
memory[2020] = 32'd5834946;
memory[2021] = 32'd7009719;
memory[2022] = 32'd6795367;
memory[2023] = 32'd8150212;
memory[2024] = 32'd5787096;
memory[2025] = 32'd833934;
memory[2026] = 32'd2019540;
memory[2027] = 32'd4221117;
memory[2028] = 32'd4726095;
memory[2029] = 32'd7278674;
memory[2030] = 32'd9473950;
memory[2031] = 32'd9520631;
memory[2032] = 32'd5728802;
memory[2033] = 32'd7727208;
memory[2034] = 32'd593630;
memory[2035] = 32'd7312851;
memory[2036] = 32'd5210525;
memory[2037] = 32'd9999242;
memory[2038] = 32'd1079690;
memory[2039] = 32'd9114447;
memory[2040] = 32'd6071161;
memory[2041] = 32'd232676;
memory[2042] = 32'd2327934;
memory[2043] = 32'd7484169;
memory[2044] = 32'd4384795;
memory[2045] = 32'd4790563;
memory[2046] = 32'd481135;
memory[2047] = 32'd5154931;
memory[2048] = 32'd9527351;
memory[2049] = 32'd776180;
memory[2050] = 32'd4541320;
memory[2051] = 32'd5362297;
memory[2052] = 32'd7785900;
memory[2053] = 32'd1336688;
memory[2054] = 32'd6028861;
memory[2055] = 32'd3572996;
memory[2056] = 32'd4686974;
memory[2057] = 32'd8048401;
memory[2058] = 32'd7794114;
memory[2059] = 32'd9413069;
memory[2060] = 32'd7843428;
memory[2061] = 32'd9784416;
memory[2062] = 32'd1450052;
memory[2063] = 32'd6088582;
memory[2064] = 32'd7511625;
memory[2065] = 32'd2043682;
memory[2066] = 32'd3401433;
memory[2067] = 32'd5238502;
memory[2068] = 32'd4559277;
memory[2069] = 32'd4481123;
memory[2070] = 32'd4352949;
memory[2071] = 32'd3146790;
memory[2072] = 32'd7230151;
memory[2073] = 32'd9197235;
memory[2074] = 32'd630960;
memory[2075] = 32'd1614946;
memory[2076] = 32'd3987799;
memory[2077] = 32'd3628447;
memory[2078] = 32'd9286229;
memory[2079] = 32'd6031502;
memory[2080] = 32'd4404628;
memory[2081] = 32'd3827549;
memory[2082] = 32'd1393799;
memory[2083] = 32'd2190528;
memory[2084] = 32'd7680589;
memory[2085] = 32'd9939013;
memory[2086] = 32'd8279876;
memory[2087] = 32'd2367563;
memory[2088] = 32'd503766;
memory[2089] = 32'd6073990;
memory[2090] = 32'd4296984;
memory[2091] = 32'd8347194;
memory[2092] = 32'd8374759;
memory[2093] = 32'd5747036;
memory[2094] = 32'd4435776;
memory[2095] = 32'd5886384;
memory[2096] = 32'd307071;
memory[2097] = 32'd7837209;
memory[2098] = 32'd3641238;
memory[2099] = 32'd7382700;
memory[2100] = 32'd4834684;
memory[2101] = 32'd510539;
memory[2102] = 32'd529490;
memory[2103] = 32'd2064835;
memory[2104] = 32'd9707775;
memory[2105] = 32'd1160450;
memory[2106] = 32'd3679781;
memory[2107] = 32'd6211926;
memory[2108] = 32'd7305250;
memory[2109] = 32'd5482362;
memory[2110] = 32'd2243428;
memory[2111] = 32'd1709878;
memory[2112] = 32'd1826264;
memory[2113] = 32'd6153579;
memory[2114] = 32'd6416758;
memory[2115] = 32'd9506853;
memory[2116] = 32'd8608944;
memory[2117] = 32'd4696634;
memory[2118] = 32'd4390769;
memory[2119] = 32'd9112711;
memory[2120] = 32'd3286977;
memory[2121] = 32'd1204105;
memory[2122] = 32'd9976257;
memory[2123] = 32'd1661736;
memory[2124] = 32'd6951142;
memory[2125] = 32'd4412034;
memory[2126] = 32'd64472;
memory[2127] = 32'd9774565;
memory[2128] = 32'd4765595;
memory[2129] = 32'd3705710;
memory[2130] = 32'd7157265;
memory[2131] = 32'd2116632;
memory[2132] = 32'd4216249;
memory[2133] = 32'd203107;
memory[2134] = 32'd4181467;
memory[2135] = 32'd6440376;
memory[2136] = 32'd1363558;
memory[2137] = 32'd377601;
memory[2138] = 32'd2652302;
memory[2139] = 32'd1185160;
memory[2140] = 32'd5859963;
memory[2141] = 32'd7412082;
memory[2142] = 32'd2895038;
memory[2143] = 32'd7686227;
memory[2144] = 32'd6082014;
memory[2145] = 32'd9311796;
memory[2146] = 32'd9709433;
memory[2147] = 32'd4690958;
memory[2148] = 32'd4008430;
memory[2149] = 32'd6616554;
memory[2150] = 32'd3803669;
memory[2151] = 32'd7295407;
memory[2152] = 32'd7820659;
memory[2153] = 32'd3779927;
memory[2154] = 32'd1473495;
memory[2155] = 32'd4771801;
memory[2156] = 32'd708313;
memory[2157] = 32'd1537967;
memory[2158] = 32'd7062718;
memory[2159] = 32'd7990260;
memory[2160] = 32'd7760029;
memory[2161] = 32'd6736335;
memory[2162] = 32'd106892;
memory[2163] = 32'd4492631;
memory[2164] = 32'd6939443;
memory[2165] = 32'd6804712;
memory[2166] = 32'd933007;
memory[2167] = 32'd819353;
memory[2168] = 32'd7182313;
memory[2169] = 32'd6101662;
memory[2170] = 32'd2004513;
memory[2171] = 32'd5558628;
memory[2172] = 32'd6030096;
memory[2173] = 32'd4899551;
memory[2174] = 32'd3244856;
memory[2175] = 32'd2112110;
memory[2176] = 32'd6727699;
memory[2177] = 32'd5470641;
memory[2178] = 32'd6803069;
memory[2179] = 32'd3252481;
memory[2180] = 32'd2087195;
memory[2181] = 32'd3123090;
memory[2182] = 32'd547889;
memory[2183] = 32'd9907854;
memory[2184] = 32'd9419369;
memory[2185] = 32'd4537736;
memory[2186] = 32'd7196008;
memory[2187] = 32'd127682;
memory[2188] = 32'd6075704;
memory[2189] = 32'd4258726;
memory[2190] = 32'd634295;
memory[2191] = 32'd3835733;
memory[2192] = 32'd3511414;
memory[2193] = 32'd741187;
memory[2194] = 32'd8328364;
memory[2195] = 32'd450857;
memory[2196] = 32'd62251;
memory[2197] = 32'd1777724;
memory[2198] = 32'd1270210;
memory[2199] = 32'd7244564;
memory[2200] = 32'd395738;
memory[2201] = 32'd3274723;
memory[2202] = 32'd2803193;
memory[2203] = 32'd6425834;
memory[2204] = 32'd690626;
memory[2205] = 32'd8564401;
memory[2206] = 32'd8537945;
memory[2207] = 32'd7418325;
memory[2208] = 32'd6551394;
memory[2209] = 32'd7857366;
memory[2210] = 32'd670806;
memory[2211] = 32'd8638589;
memory[2212] = 32'd980456;
memory[2213] = 32'd3735047;
memory[2214] = 32'd1062795;
memory[2215] = 32'd399826;
memory[2216] = 32'd8272784;
memory[2217] = 32'd8258803;
memory[2218] = 32'd3043860;
memory[2219] = 32'd6864840;
memory[2220] = 32'd5033882;
memory[2221] = 32'd3678155;
memory[2222] = 32'd700573;
memory[2223] = 32'd1061648;
memory[2224] = 32'd6935695;
memory[2225] = 32'd1545290;
memory[2226] = 32'd1512505;
memory[2227] = 32'd6997946;
memory[2228] = 32'd5839366;
memory[2229] = 32'd5299067;
memory[2230] = 32'd6758863;
memory[2231] = 32'd6235104;
memory[2232] = 32'd8573790;
memory[2233] = 32'd2078408;
memory[2234] = 32'd5177290;
memory[2235] = 32'd1780768;
memory[2236] = 32'd3159161;
memory[2237] = 32'd3715235;
memory[2238] = 32'd9199093;
memory[2239] = 32'd9710555;
memory[2240] = 32'd1572601;
memory[2241] = 32'd2386251;
memory[2242] = 32'd8349144;
memory[2243] = 32'd5069410;
memory[2244] = 32'd8637651;
memory[2245] = 32'd1928291;
memory[2246] = 32'd7985588;
memory[2247] = 32'd6910435;
memory[2248] = 32'd2703447;
memory[2249] = 32'd1029448;
memory[2250] = 32'd3775275;
memory[2251] = 32'd253681;
memory[2252] = 32'd7223956;
memory[2253] = 32'd6992200;
memory[2254] = 32'd1315329;
memory[2255] = 32'd4159651;
memory[2256] = 32'd1053842;
memory[2257] = 32'd2827834;
memory[2258] = 32'd3673949;
memory[2259] = 32'd9409560;
memory[2260] = 32'd8126901;
memory[2261] = 32'd2949164;
memory[2262] = 32'd5644664;
memory[2263] = 32'd9217043;
memory[2264] = 32'd5027572;
memory[2265] = 32'd821955;
memory[2266] = 32'd997811;
memory[2267] = 32'd8186733;
memory[2268] = 32'd7053542;
memory[2269] = 32'd2713256;
memory[2270] = 32'd413640;
memory[2271] = 32'd1142496;
memory[2272] = 32'd7615859;
memory[2273] = 32'd1279136;
memory[2274] = 32'd8728258;
memory[2275] = 32'd6253510;
memory[2276] = 32'd3207428;
memory[2277] = 32'd6713846;
memory[2278] = 32'd5680297;
memory[2279] = 32'd5910875;
memory[2280] = 32'd7743294;
memory[2281] = 32'd1971924;
memory[2282] = 32'd6164556;
memory[2283] = 32'd4967250;
memory[2284] = 32'd8964125;
memory[2285] = 32'd7479885;
memory[2286] = 32'd1643253;
memory[2287] = 32'd2534319;
memory[2288] = 32'd2824071;
memory[2289] = 32'd7833555;
memory[2290] = 32'd1943880;
memory[2291] = 32'd3467324;
memory[2292] = 32'd782719;
memory[2293] = 32'd104896;
memory[2294] = 32'd2684367;
memory[2295] = 32'd8326644;
memory[2296] = 32'd3443203;
memory[2297] = 32'd6198530;
memory[2298] = 32'd9029729;
memory[2299] = 32'd496746;
memory[2300] = 32'd8911786;
memory[2301] = 32'd9443370;
memory[2302] = 32'd4155594;
memory[2303] = 32'd6527645;
memory[2304] = 32'd3238858;
memory[2305] = 32'd2883852;
memory[2306] = 32'd5297508;
memory[2307] = 32'd6446286;
memory[2308] = 32'd9597698;
memory[2309] = 32'd977805;
memory[2310] = 32'd4873513;
memory[2311] = 32'd9857344;
memory[2312] = 32'd2949730;
memory[2313] = 32'd3554421;
memory[2314] = 32'd7340947;
memory[2315] = 32'd4430207;
memory[2316] = 32'd3550658;
memory[2317] = 32'd8984200;
memory[2318] = 32'd9480878;
memory[2319] = 32'd6374729;
memory[2320] = 32'd9334107;
memory[2321] = 32'd1424758;
memory[2322] = 32'd9842053;
memory[2323] = 32'd2633179;
memory[2324] = 32'd4046007;
memory[2325] = 32'd5042772;
memory[2326] = 32'd3476175;
memory[2327] = 32'd7489210;
memory[2328] = 32'd1241302;
memory[2329] = 32'd2505904;
memory[2330] = 32'd502308;
memory[2331] = 32'd2669440;
memory[2332] = 32'd4465626;
memory[2333] = 32'd4657902;
memory[2334] = 32'd9197086;
memory[2335] = 32'd7704485;
memory[2336] = 32'd58106;
memory[2337] = 32'd7010946;
memory[2338] = 32'd6667123;
memory[2339] = 32'd9655804;
memory[2340] = 32'd7988751;
memory[2341] = 32'd1540637;
memory[2342] = 32'd2029501;
memory[2343] = 32'd3454833;
memory[2344] = 32'd7611410;
memory[2345] = 32'd9370448;
memory[2346] = 32'd401392;
memory[2347] = 32'd1162069;
memory[2348] = 32'd871000;
memory[2349] = 32'd9882271;
memory[2350] = 32'd53150;
memory[2351] = 32'd205108;
memory[2352] = 32'd3823381;
memory[2353] = 32'd2411556;
memory[2354] = 32'd2838287;
memory[2355] = 32'd7869388;
memory[2356] = 32'd7454328;
memory[2357] = 32'd6314462;
memory[2358] = 32'd7874951;
memory[2359] = 32'd1211983;
memory[2360] = 32'd1336718;
memory[2361] = 32'd8377259;
memory[2362] = 32'd3881423;
memory[2363] = 32'd5802345;
memory[2364] = 32'd5551514;
memory[2365] = 32'd5594861;
memory[2366] = 32'd6023182;
memory[2367] = 32'd8125972;
memory[2368] = 32'd2605807;
memory[2369] = 32'd5206657;
memory[2370] = 32'd298129;
memory[2371] = 32'd3110911;
memory[2372] = 32'd6747294;
memory[2373] = 32'd2327630;
memory[2374] = 32'd6565744;
memory[2375] = 32'd6875057;
memory[2376] = 32'd1698078;
memory[2377] = 32'd6967137;
memory[2378] = 32'd8037126;
memory[2379] = 32'd2569078;
memory[2380] = 32'd9365760;
memory[2381] = 32'd606628;
memory[2382] = 32'd2774186;
memory[2383] = 32'd3189141;
memory[2384] = 32'd3018184;
memory[2385] = 32'd8128825;
memory[2386] = 32'd3574882;
memory[2387] = 32'd2988865;
memory[2388] = 32'd6959639;
memory[2389] = 32'd1449833;
memory[2390] = 32'd4200848;
memory[2391] = 32'd8296358;
memory[2392] = 32'd2343444;
memory[2393] = 32'd598623;
memory[2394] = 32'd6615055;
memory[2395] = 32'd411310;
memory[2396] = 32'd6193485;
memory[2397] = 32'd5154589;
memory[2398] = 32'd8537283;
memory[2399] = 32'd1315644;
memory[2400] = 32'd361246;
memory[2401] = 32'd8835412;
memory[2402] = 32'd4426555;
memory[2403] = 32'd9624893;
memory[2404] = 32'd1163042;
memory[2405] = 32'd992300;
memory[2406] = 32'd6499950;
memory[2407] = 32'd2861120;
memory[2408] = 32'd475789;
memory[2409] = 32'd7053428;
memory[2410] = 32'd7946550;
memory[2411] = 32'd9841549;
memory[2412] = 32'd7660056;
memory[2413] = 32'd720737;
memory[2414] = 32'd5547042;
memory[2415] = 32'd678241;
memory[2416] = 32'd1365914;
memory[2417] = 32'd9121924;
memory[2418] = 32'd6183458;
memory[2419] = 32'd8325554;
memory[2420] = 32'd3088109;
memory[2421] = 32'd2900658;
memory[2422] = 32'd9138264;
memory[2423] = 32'd5431554;
memory[2424] = 32'd3499281;
memory[2425] = 32'd5753319;
memory[2426] = 32'd8359216;
memory[2427] = 32'd2209118;
memory[2428] = 32'd3424260;
memory[2429] = 32'd6896499;
memory[2430] = 32'd3524763;
memory[2431] = 32'd3785506;
memory[2432] = 32'd8248263;
memory[2433] = 32'd7951318;
memory[2434] = 32'd3410399;
memory[2435] = 32'd9411305;
memory[2436] = 32'd1459970;
memory[2437] = 32'd2426701;
memory[2438] = 32'd4788777;
memory[2439] = 32'd4452111;
memory[2440] = 32'd9480129;
memory[2441] = 32'd2735328;
memory[2442] = 32'd6810012;
memory[2443] = 32'd7140186;
memory[2444] = 32'd5972417;
memory[2445] = 32'd2357055;
memory[2446] = 32'd334779;
memory[2447] = 32'd9854683;
memory[2448] = 32'd1478979;
memory[2449] = 32'd9034589;
memory[2450] = 32'd8180237;
memory[2451] = 32'd4567089;
memory[2452] = 32'd1935247;
memory[2453] = 32'd9834853;
memory[2454] = 32'd2514995;
memory[2455] = 32'd7950880;
memory[2456] = 32'd8104524;
memory[2457] = 32'd874211;
memory[2458] = 32'd159999;
memory[2459] = 32'd1528784;
memory[2460] = 32'd7770711;
memory[2461] = 32'd6201114;
memory[2462] = 32'd7830643;
memory[2463] = 32'd8535326;
memory[2464] = 32'd6668784;
memory[2465] = 32'd1241042;
memory[2466] = 32'd7946632;
memory[2467] = 32'd645107;
memory[2468] = 32'd6184096;
memory[2469] = 32'd5251761;
memory[2470] = 32'd5097218;
memory[2471] = 32'd5664225;
memory[2472] = 32'd503441;
memory[2473] = 32'd1907231;
memory[2474] = 32'd5320763;
memory[2475] = 32'd8992210;
memory[2476] = 32'd4264286;
memory[2477] = 32'd8171894;
memory[2478] = 32'd8846894;
memory[2479] = 32'd8259617;
memory[2480] = 32'd9722835;
memory[2481] = 32'd9543483;
memory[2482] = 32'd5343058;
memory[2483] = 32'd1658082;
memory[2484] = 32'd9378337;
memory[2485] = 32'd7858053;
memory[2486] = 32'd2125315;
memory[2487] = 32'd9999213;
memory[2488] = 32'd1248617;
memory[2489] = 32'd2285314;
memory[2490] = 32'd1527998;
memory[2491] = 32'd1535680;
memory[2492] = 32'd1002780;
memory[2493] = 32'd9358641;
memory[2494] = 32'd71006;
memory[2495] = 32'd7671564;
memory[2496] = 32'd3116035;
memory[2497] = 32'd8017638;
memory[2498] = 32'd833023;
memory[2499] = 32'd9300131;
memory[2500] = 32'd5785752;
memory[2501] = 32'd5930242;
memory[2502] = 32'd7480709;
memory[2503] = 32'd8805545;
memory[2504] = 32'd353825;
memory[2505] = 32'd5317824;
memory[2506] = 32'd7797756;
memory[2507] = 32'd7134463;
memory[2508] = 32'd6006071;
memory[2509] = 32'd9161002;
memory[2510] = 32'd5394080;
memory[2511] = 32'd5728906;
memory[2512] = 32'd8704485;
memory[2513] = 32'd3253491;
memory[2514] = 32'd7386989;
memory[2515] = 32'd599174;
memory[2516] = 32'd1111544;
memory[2517] = 32'd2028656;
memory[2518] = 32'd598388;
memory[2519] = 32'd2360161;
memory[2520] = 32'd4313970;
memory[2521] = 32'd4642738;
memory[2522] = 32'd3895841;
memory[2523] = 32'd7833102;
memory[2524] = 32'd4001379;
memory[2525] = 32'd3966848;
memory[2526] = 32'd8021018;
memory[2527] = 32'd9633766;
memory[2528] = 32'd4500838;
memory[2529] = 32'd8854042;
memory[2530] = 32'd1450250;
memory[2531] = 32'd2802942;
memory[2532] = 32'd4784284;
memory[2533] = 32'd8930959;
memory[2534] = 32'd1608488;
memory[2535] = 32'd7654461;
memory[2536] = 32'd6765135;
memory[2537] = 32'd1922596;
memory[2538] = 32'd4788924;
memory[2539] = 32'd2771206;
memory[2540] = 32'd1083598;
memory[2541] = 32'd2699356;
memory[2542] = 32'd8500113;
memory[2543] = 32'd2304435;
memory[2544] = 32'd5952847;
memory[2545] = 32'd8403454;
memory[2546] = 32'd5419962;
memory[2547] = 32'd9580744;
memory[2548] = 32'd432110;
memory[2549] = 32'd8534702;
memory[2550] = 32'd4457257;
memory[2551] = 32'd7262432;
memory[2552] = 32'd3177440;
memory[2553] = 32'd869451;
memory[2554] = 32'd7611886;
memory[2555] = 32'd9695171;
memory[2556] = 32'd4836299;
memory[2557] = 32'd5632904;
memory[2558] = 32'd1845289;
memory[2559] = 32'd1853489;
memory[2560] = 32'd4486946;
memory[2561] = 32'd3295539;
memory[2562] = 32'd7172784;
memory[2563] = 32'd1787582;
memory[2564] = 32'd4742850;
memory[2565] = 32'd8781272;
memory[2566] = 32'd9442043;
memory[2567] = 32'd1507986;
memory[2568] = 32'd703868;
memory[2569] = 32'd6747319;
memory[2570] = 32'd4279192;
memory[2571] = 32'd4303818;
memory[2572] = 32'd9446676;
memory[2573] = 32'd5295657;
memory[2574] = 32'd6608253;
memory[2575] = 32'd7915875;
memory[2576] = 32'd6215463;
memory[2577] = 32'd2028215;
memory[2578] = 32'd7496619;
memory[2579] = 32'd9163925;
memory[2580] = 32'd3079269;
memory[2581] = 32'd1953877;
memory[2582] = 32'd8942709;
memory[2583] = 32'd6256709;
memory[2584] = 32'd5339680;
memory[2585] = 32'd6554595;
memory[2586] = 32'd8468232;
memory[2587] = 32'd2692331;
memory[2588] = 32'd2187500;
memory[2589] = 32'd313522;
memory[2590] = 32'd4545820;
memory[2591] = 32'd6674446;
memory[2592] = 32'd6125413;
memory[2593] = 32'd4234956;
memory[2594] = 32'd8462029;
memory[2595] = 32'd868264;
memory[2596] = 32'd3016228;
memory[2597] = 32'd420424;
memory[2598] = 32'd2376250;
memory[2599] = 32'd6236448;
memory[2600] = 32'd7167744;
memory[2601] = 32'd9171794;
memory[2602] = 32'd3056618;
memory[2603] = 32'd9130772;
memory[2604] = 32'd6983804;
memory[2605] = 32'd9664872;
memory[2606] = 32'd7046647;
memory[2607] = 32'd3199267;
memory[2608] = 32'd4209439;
memory[2609] = 32'd7059619;
memory[2610] = 32'd2363193;
memory[2611] = 32'd7288709;
memory[2612] = 32'd1529848;
memory[2613] = 32'd3822254;
memory[2614] = 32'd6061770;
memory[2615] = 32'd6869528;
memory[2616] = 32'd376850;
memory[2617] = 32'd7046355;
memory[2618] = 32'd9561859;
memory[2619] = 32'd2564350;
memory[2620] = 32'd9876229;
memory[2621] = 32'd6624031;
memory[2622] = 32'd1755148;
memory[2623] = 32'd6001642;
memory[2624] = 32'd858988;
memory[2625] = 32'd217177;
memory[2626] = 32'd6869906;
memory[2627] = 32'd6391568;
memory[2628] = 32'd3153954;
memory[2629] = 32'd1762508;
memory[2630] = 32'd5144369;
memory[2631] = 32'd321698;
memory[2632] = 32'd934303;
memory[2633] = 32'd8200987;
memory[2634] = 32'd9452470;
memory[2635] = 32'd7918107;
memory[2636] = 32'd382211;
memory[2637] = 32'd9015469;
memory[2638] = 32'd3633726;
memory[2639] = 32'd7108003;
memory[2640] = 32'd8591440;
memory[2641] = 32'd8513271;
memory[2642] = 32'd6913064;
memory[2643] = 32'd121288;
memory[2644] = 32'd2335526;
memory[2645] = 32'd5491186;
memory[2646] = 32'd6990816;
memory[2647] = 32'd2712376;
memory[2648] = 32'd2537541;
memory[2649] = 32'd9069027;
memory[2650] = 32'd7793078;
memory[2651] = 32'd4930122;
memory[2652] = 32'd5693059;
memory[2653] = 32'd9548226;
memory[2654] = 32'd931765;
memory[2655] = 32'd9068399;
memory[2656] = 32'd9765404;
memory[2657] = 32'd318023;
memory[2658] = 32'd5459967;
memory[2659] = 32'd2919358;
memory[2660] = 32'd2080532;
memory[2661] = 32'd3120688;
memory[2662] = 32'd5757408;
memory[2663] = 32'd5531187;
memory[2664] = 32'd1321676;
memory[2665] = 32'd7726230;
memory[2666] = 32'd3449294;
memory[2667] = 32'd4220239;
memory[2668] = 32'd9258051;
memory[2669] = 32'd9599372;
memory[2670] = 32'd1328242;
memory[2671] = 32'd7849492;
memory[2672] = 32'd8112644;
memory[2673] = 32'd8241306;
memory[2674] = 32'd7970780;
memory[2675] = 32'd2964522;
memory[2676] = 32'd3732493;
memory[2677] = 32'd7477949;
memory[2678] = 32'd5676898;
memory[2679] = 32'd8786386;
memory[2680] = 32'd9063328;
memory[2681] = 32'd3469976;
memory[2682] = 32'd3716509;
memory[2683] = 32'd4756387;
memory[2684] = 32'd3018202;
memory[2685] = 32'd7164626;
memory[2686] = 32'd6341138;
memory[2687] = 32'd5299958;
memory[2688] = 32'd7482649;
memory[2689] = 32'd4317458;
memory[2690] = 32'd735668;
memory[2691] = 32'd9563181;
memory[2692] = 32'd7438146;
memory[2693] = 32'd9009428;
memory[2694] = 32'd7610720;
memory[2695] = 32'd1276174;
memory[2696] = 32'd6735658;
memory[2697] = 32'd1060014;
memory[2698] = 32'd5496414;
memory[2699] = 32'd8510062;
memory[2700] = 32'd3175739;
memory[2701] = 32'd6824656;
memory[2702] = 32'd6359554;
memory[2703] = 32'd3804735;
memory[2704] = 32'd7582315;
memory[2705] = 32'd4330334;
memory[2706] = 32'd6769257;
memory[2707] = 32'd3831160;
memory[2708] = 32'd4324635;
memory[2709] = 32'd4962507;
memory[2710] = 32'd2617546;
memory[2711] = 32'd3387964;
memory[2712] = 32'd8432483;
memory[2713] = 32'd6334055;
memory[2714] = 32'd660703;
memory[2715] = 32'd3967037;
memory[2716] = 32'd6015033;
memory[2717] = 32'd7001842;
memory[2718] = 32'd1783348;
memory[2719] = 32'd3497683;
memory[2720] = 32'd1319300;
memory[2721] = 32'd5035368;
memory[2722] = 32'd5577216;
memory[2723] = 32'd8757446;
memory[2724] = 32'd6561149;
memory[2725] = 32'd3187937;
memory[2726] = 32'd33621;
memory[2727] = 32'd5813159;
memory[2728] = 32'd6764303;
memory[2729] = 32'd8046387;
memory[2730] = 32'd4323221;
memory[2731] = 32'd9940042;
memory[2732] = 32'd4871043;
memory[2733] = 32'd682775;
memory[2734] = 32'd3744777;
memory[2735] = 32'd4969710;
memory[2736] = 32'd7529462;
memory[2737] = 32'd3030386;
memory[2738] = 32'd8800870;
memory[2739] = 32'd1854097;
memory[2740] = 32'd7992893;
memory[2741] = 32'd1418417;
memory[2742] = 32'd5242061;
memory[2743] = 32'd8941728;
memory[2744] = 32'd268824;
memory[2745] = 32'd8419117;
memory[2746] = 32'd2908766;
memory[2747] = 32'd6283858;
memory[2748] = 32'd5420959;
memory[2749] = 32'd7208466;
memory[2750] = 32'd2297893;
memory[2751] = 32'd6740259;
memory[2752] = 32'd4760186;
memory[2753] = 32'd7875109;
memory[2754] = 32'd8014057;
memory[2755] = 32'd1321335;
memory[2756] = 32'd1063046;
memory[2757] = 32'd564030;
memory[2758] = 32'd7134495;
memory[2759] = 32'd343702;
memory[2760] = 32'd8610417;
memory[2761] = 32'd1457716;
memory[2762] = 32'd2800096;
memory[2763] = 32'd5997813;
memory[2764] = 32'd2140492;
memory[2765] = 32'd6544874;
memory[2766] = 32'd967523;
memory[2767] = 32'd2186306;
memory[2768] = 32'd9575260;
memory[2769] = 32'd9768394;
memory[2770] = 32'd4040403;
memory[2771] = 32'd84506;
memory[2772] = 32'd3703163;
memory[2773] = 32'd1798817;
memory[2774] = 32'd9026234;
memory[2775] = 32'd6488339;
memory[2776] = 32'd217934;
memory[2777] = 32'd4451352;
memory[2778] = 32'd5288549;
memory[2779] = 32'd5638893;
memory[2780] = 32'd1659818;
memory[2781] = 32'd7586442;
memory[2782] = 32'd4895504;
memory[2783] = 32'd6420005;
memory[2784] = 32'd7977904;
memory[2785] = 32'd5425913;
memory[2786] = 32'd257692;
memory[2787] = 32'd1557302;
memory[2788] = 32'd5989944;
memory[2789] = 32'd7392187;
memory[2790] = 32'd1901004;
memory[2791] = 32'd4600361;
memory[2792] = 32'd1366256;
memory[2793] = 32'd4701101;
memory[2794] = 32'd3114526;
memory[2795] = 32'd3506748;
memory[2796] = 32'd3762327;
memory[2797] = 32'd4082050;
memory[2798] = 32'd5693054;
memory[2799] = 32'd5853939;
memory[2800] = 32'd6366796;
memory[2801] = 32'd2249809;
memory[2802] = 32'd5938445;
memory[2803] = 32'd2586311;
memory[2804] = 32'd4048626;
memory[2805] = 32'd4964680;
memory[2806] = 32'd1591002;
memory[2807] = 32'd6782912;
memory[2808] = 32'd9416032;
memory[2809] = 32'd6879552;
memory[2810] = 32'd4938157;
memory[2811] = 32'd3592203;
memory[2812] = 32'd6982346;
memory[2813] = 32'd9833661;
memory[2814] = 32'd2528560;
memory[2815] = 32'd4960250;
memory[2816] = 32'd7775927;
memory[2817] = 32'd2786252;
memory[2818] = 32'd6517553;
memory[2819] = 32'd3765871;
memory[2820] = 32'd178440;
memory[2821] = 32'd8418557;
memory[2822] = 32'd882584;
memory[2823] = 32'd4061048;
memory[2824] = 32'd5636010;
memory[2825] = 32'd3997111;
memory[2826] = 32'd84148;
memory[2827] = 32'd9398337;
memory[2828] = 32'd595513;
memory[2829] = 32'd8293554;
memory[2830] = 32'd5252277;
memory[2831] = 32'd9478661;
memory[2832] = 32'd543363;
memory[2833] = 32'd3707074;
memory[2834] = 32'd4581324;
memory[2835] = 32'd7108342;
memory[2836] = 32'd8671754;
memory[2837] = 32'd6172326;
memory[2838] = 32'd3891254;
memory[2839] = 32'd604139;
memory[2840] = 32'd3051878;
memory[2841] = 32'd1345764;
memory[2842] = 32'd4196342;
memory[2843] = 32'd34225;
memory[2844] = 32'd3695777;
memory[2845] = 32'd6724902;
memory[2846] = 32'd7510827;
memory[2847] = 32'd1471704;
memory[2848] = 32'd9511154;
memory[2849] = 32'd4028380;
memory[2850] = 32'd5237575;
memory[2851] = 32'd2205946;
memory[2852] = 32'd4963290;
memory[2853] = 32'd6120160;
memory[2854] = 32'd6266994;
memory[2855] = 32'd599300;
memory[2856] = 32'd2633623;
memory[2857] = 32'd6351142;
memory[2858] = 32'd2513990;
memory[2859] = 32'd5745488;
memory[2860] = 32'd4644696;
memory[2861] = 32'd282619;
memory[2862] = 32'd5224149;
memory[2863] = 32'd7704412;
memory[2864] = 32'd3989693;
memory[2865] = 32'd2321825;
memory[2866] = 32'd4812754;
memory[2867] = 32'd2661448;
memory[2868] = 32'd8494151;
memory[2869] = 32'd1220360;
memory[2870] = 32'd3265587;
memory[2871] = 32'd4062382;
memory[2872] = 32'd2566124;
memory[2873] = 32'd7461929;
memory[2874] = 32'd6612959;
memory[2875] = 32'd6261902;
memory[2876] = 32'd6703183;
memory[2877] = 32'd4123786;
memory[2878] = 32'd7733606;
memory[2879] = 32'd6214337;
memory[2880] = 32'd8152167;
memory[2881] = 32'd5487534;
memory[2882] = 32'd936636;
memory[2883] = 32'd5631809;
memory[2884] = 32'd4124046;
memory[2885] = 32'd7203630;
memory[2886] = 32'd6231109;
memory[2887] = 32'd6757669;
memory[2888] = 32'd6071125;
memory[2889] = 32'd1261451;
memory[2890] = 32'd2503157;
memory[2891] = 32'd3232173;
memory[2892] = 32'd1544070;
memory[2893] = 32'd243658;
memory[2894] = 32'd936585;
memory[2895] = 32'd5533764;
memory[2896] = 32'd2565483;
memory[2897] = 32'd5749339;
memory[2898] = 32'd711564;
memory[2899] = 32'd3575986;
memory[2900] = 32'd9486052;
memory[2901] = 32'd6493503;
memory[2902] = 32'd7638368;
memory[2903] = 32'd2052176;
memory[2904] = 32'd3955432;
memory[2905] = 32'd4251327;
memory[2906] = 32'd830430;
memory[2907] = 32'd3174967;
memory[2908] = 32'd891466;
memory[2909] = 32'd8564037;
memory[2910] = 32'd9389304;
memory[2911] = 32'd9043633;
memory[2912] = 32'd4051571;
memory[2913] = 32'd2842292;
memory[2914] = 32'd7191794;
memory[2915] = 32'd8175617;
memory[2916] = 32'd2562275;
memory[2917] = 32'd5939255;
memory[2918] = 32'd7449638;
memory[2919] = 32'd8633400;
memory[2920] = 32'd7200707;
memory[2921] = 32'd2469147;
memory[2922] = 32'd1865573;
memory[2923] = 32'd8744777;
memory[2924] = 32'd5229157;
memory[2925] = 32'd2802159;
memory[2926] = 32'd6794893;
memory[2927] = 32'd310992;
memory[2928] = 32'd1067850;
memory[2929] = 32'd7506457;
memory[2930] = 32'd3886978;
memory[2931] = 32'd553902;
memory[2932] = 32'd3999960;
memory[2933] = 32'd1525347;
memory[2934] = 32'd5122431;
memory[2935] = 32'd471744;
memory[2936] = 32'd8293026;
memory[2937] = 32'd5952861;
memory[2938] = 32'd3646711;
memory[2939] = 32'd9184492;
memory[2940] = 32'd4516898;
memory[2941] = 32'd5552368;
memory[2942] = 32'd744477;
memory[2943] = 32'd1084821;
memory[2944] = 32'd8394660;
memory[2945] = 32'd7936271;
memory[2946] = 32'd1776790;
memory[2947] = 32'd3473287;
memory[2948] = 32'd6391879;
memory[2949] = 32'd1742780;
memory[2950] = 32'd2106687;
memory[2951] = 32'd3592586;
memory[2952] = 32'd6728279;
memory[2953] = 32'd6488613;
memory[2954] = 32'd2337363;
memory[2955] = 32'd1957436;
memory[2956] = 32'd1807124;
memory[2957] = 32'd1648609;
memory[2958] = 32'd2268428;
memory[2959] = 32'd2874974;
memory[2960] = 32'd9155066;
memory[2961] = 32'd8671759;
memory[2962] = 32'd5945229;
memory[2963] = 32'd3155027;
memory[2964] = 32'd2713458;
memory[2965] = 32'd1067660;
memory[2966] = 32'd3626771;
memory[2967] = 32'd1006484;
memory[2968] = 32'd9536873;
memory[2969] = 32'd9789835;
memory[2970] = 32'd2707329;
memory[2971] = 32'd6570124;
memory[2972] = 32'd5342203;
memory[2973] = 32'd5968158;
memory[2974] = 32'd7654945;
memory[2975] = 32'd6253215;
memory[2976] = 32'd6420782;
memory[2977] = 32'd1948088;
memory[2978] = 32'd9726503;
memory[2979] = 32'd2812661;
memory[2980] = 32'd3690868;
memory[2981] = 32'd4349542;
memory[2982] = 32'd6405247;
memory[2983] = 32'd2935500;
memory[2984] = 32'd838155;
memory[2985] = 32'd1258962;
memory[2986] = 32'd4892936;
memory[2987] = 32'd5161631;
memory[2988] = 32'd2907571;
memory[2989] = 32'd9677717;
memory[2990] = 32'd552958;
memory[2991] = 32'd2062638;
memory[2992] = 32'd8349476;
memory[2993] = 32'd6498187;
memory[2994] = 32'd7734017;
memory[2995] = 32'd1062934;
memory[2996] = 32'd82199;
memory[2997] = 32'd3877140;
memory[2998] = 32'd4585770;
memory[2999] = 32'd9619072;
memory[3000] = 32'd6183327;
memory[3001] = 32'd9809451;
memory[3002] = 32'd6189196;
memory[3003] = 32'd4041882;
memory[3004] = 32'd5777610;
memory[3005] = 32'd6360494;
memory[3006] = 32'd295098;
memory[3007] = 32'd2198392;
memory[3008] = 32'd8308582;
memory[3009] = 32'd2537953;
memory[3010] = 32'd5011053;
memory[3011] = 32'd4515802;
memory[3012] = 32'd9403847;
memory[3013] = 32'd3932652;
memory[3014] = 32'd9967654;
memory[3015] = 32'd2758355;
memory[3016] = 32'd5191614;
memory[3017] = 32'd4860591;
memory[3018] = 32'd7919986;
memory[3019] = 32'd615538;
memory[3020] = 32'd7054660;
memory[3021] = 32'd8472944;
memory[3022] = 32'd5194528;
memory[3023] = 32'd7920488;
memory[3024] = 32'd7487483;
memory[3025] = 32'd2928545;
memory[3026] = 32'd8983422;
memory[3027] = 32'd86034;
memory[3028] = 32'd9322037;
memory[3029] = 32'd6085544;
memory[3030] = 32'd9705107;
memory[3031] = 32'd5505365;
memory[3032] = 32'd5894996;
memory[3033] = 32'd8410655;
memory[3034] = 32'd9547247;
memory[3035] = 32'd1672606;
memory[3036] = 32'd4771149;
memory[3037] = 32'd2358697;
memory[3038] = 32'd6387350;
memory[3039] = 32'd5596083;
memory[3040] = 32'd7413002;
memory[3041] = 32'd1398403;
memory[3042] = 32'd2628238;
memory[3043] = 32'd6816850;
memory[3044] = 32'd5331055;
memory[3045] = 32'd2595892;
memory[3046] = 32'd9575205;
memory[3047] = 32'd3039021;
memory[3048] = 32'd9972835;
memory[3049] = 32'd7495191;
memory[3050] = 32'd6170911;
memory[3051] = 32'd7027495;
memory[3052] = 32'd8484488;
memory[3053] = 32'd1365439;
memory[3054] = 32'd4947983;
memory[3055] = 32'd8488323;
memory[3056] = 32'd6810336;
memory[3057] = 32'd6447757;
memory[3058] = 32'd8574358;
memory[3059] = 32'd8648726;
memory[3060] = 32'd2533302;
memory[3061] = 32'd8279465;
memory[3062] = 32'd4154091;
memory[3063] = 32'd944650;
memory[3064] = 32'd6690120;
memory[3065] = 32'd6217690;
memory[3066] = 32'd5133608;
memory[3067] = 32'd3977622;
memory[3068] = 32'd8576388;
memory[3069] = 32'd1520958;
memory[3070] = 32'd2090057;
memory[3071] = 32'd5989390;
memory[3072] = 32'd2919361;
memory[3073] = 32'd4718295;
memory[3074] = 32'd2806240;
memory[3075] = 32'd766768;
memory[3076] = 32'd9830540;
memory[3077] = 32'd4897797;
memory[3078] = 32'd6322141;
memory[3079] = 32'd9803375;
memory[3080] = 32'd4909341;
memory[3081] = 32'd2493053;
memory[3082] = 32'd9347223;
memory[3083] = 32'd3393829;
memory[3084] = 32'd6374844;
memory[3085] = 32'd6811558;
memory[3086] = 32'd1882152;
memory[3087] = 32'd5701533;
memory[3088] = 32'd3259316;
memory[3089] = 32'd456510;
memory[3090] = 32'd4350259;
memory[3091] = 32'd8308970;
memory[3092] = 32'd1252327;
memory[3093] = 32'd8504350;
memory[3094] = 32'd1769972;
memory[3095] = 32'd458800;
memory[3096] = 32'd4722040;
memory[3097] = 32'd6903580;
memory[3098] = 32'd6952774;
memory[3099] = 32'd5814780;
memory[3100] = 32'd8424538;
memory[3101] = 32'd9042831;
memory[3102] = 32'd1804171;
memory[3103] = 32'd1343899;
memory[3104] = 32'd6277479;
memory[3105] = 32'd7126763;
memory[3106] = 32'd4627019;
memory[3107] = 32'd6108019;
memory[3108] = 32'd2024561;
memory[3109] = 32'd3465512;
memory[3110] = 32'd8427746;
memory[3111] = 32'd9450254;
memory[3112] = 32'd8474917;
memory[3113] = 32'd7774969;
memory[3114] = 32'd2844083;
memory[3115] = 32'd4849762;
memory[3116] = 32'd4586528;
memory[3117] = 32'd7242587;
memory[3118] = 32'd551295;
memory[3119] = 32'd362196;
memory[3120] = 32'd215450;
memory[3121] = 32'd4901554;
memory[3122] = 32'd8671166;
memory[3123] = 32'd3984129;
memory[3124] = 32'd5922256;
memory[3125] = 32'd441138;
memory[3126] = 32'd4442929;
memory[3127] = 32'd644296;
memory[3128] = 32'd7344718;
memory[3129] = 32'd3912055;
memory[3130] = 32'd8975429;
memory[3131] = 32'd8285608;
memory[3132] = 32'd2954887;
memory[3133] = 32'd779600;
memory[3134] = 32'd9629507;
memory[3135] = 32'd1748718;
memory[3136] = 32'd422715;
memory[3137] = 32'd6772878;
memory[3138] = 32'd7856737;
memory[3139] = 32'd4963628;
memory[3140] = 32'd238390;
memory[3141] = 32'd8800835;
memory[3142] = 32'd4413882;
memory[3143] = 32'd8713308;
memory[3144] = 32'd6575805;
memory[3145] = 32'd9774317;
memory[3146] = 32'd6079422;
memory[3147] = 32'd3678685;
memory[3148] = 32'd9533257;
memory[3149] = 32'd9147069;
memory[3150] = 32'd4040881;
memory[3151] = 32'd9748707;
memory[3152] = 32'd4048623;
memory[3153] = 32'd5228399;
memory[3154] = 32'd3732836;
memory[3155] = 32'd9970879;
memory[3156] = 32'd8185889;
memory[3157] = 32'd692118;
memory[3158] = 32'd3131527;
memory[3159] = 32'd5530607;
memory[3160] = 32'd4604173;
memory[3161] = 32'd2106956;
memory[3162] = 32'd3816215;
memory[3163] = 32'd75412;
memory[3164] = 32'd5402908;
memory[3165] = 32'd5962074;
memory[3166] = 32'd1824130;
memory[3167] = 32'd8341976;
memory[3168] = 32'd5251304;
memory[3169] = 32'd2197219;
memory[3170] = 32'd5821956;
memory[3171] = 32'd8006046;
memory[3172] = 32'd998055;
memory[3173] = 32'd235839;
memory[3174] = 32'd9235706;
memory[3175] = 32'd90212;
memory[3176] = 32'd2526508;
memory[3177] = 32'd5315128;
memory[3178] = 32'd3768897;
memory[3179] = 32'd2059765;
memory[3180] = 32'd4462197;
memory[3181] = 32'd326130;
memory[3182] = 32'd1808472;
memory[3183] = 32'd1027172;
memory[3184] = 32'd5554529;
memory[3185] = 32'd8057661;
memory[3186] = 32'd3514403;
memory[3187] = 32'd3740418;
memory[3188] = 32'd1266131;
memory[3189] = 32'd9162283;
memory[3190] = 32'd1787377;
memory[3191] = 32'd8386656;
memory[3192] = 32'd3785591;
memory[3193] = 32'd8119944;
memory[3194] = 32'd8462069;
memory[3195] = 32'd1704852;
memory[3196] = 32'd6598370;
memory[3197] = 32'd2802551;
memory[3198] = 32'd46828;
memory[3199] = 32'd4366026;
memory[3200] = 32'd7516123;
memory[3201] = 32'd5868784;
memory[3202] = 32'd2372072;
memory[3203] = 32'd1030530;
memory[3204] = 32'd8620975;
memory[3205] = 32'd1607779;
memory[3206] = 32'd3637094;
memory[3207] = 32'd1147484;
memory[3208] = 32'd9439259;
memory[3209] = 32'd7405991;
memory[3210] = 32'd3207249;
memory[3211] = 32'd6417809;
memory[3212] = 32'd248473;
memory[3213] = 32'd7532074;
memory[3214] = 32'd7444981;
memory[3215] = 32'd5803002;
memory[3216] = 32'd5589735;
memory[3217] = 32'd3475737;
memory[3218] = 32'd2059772;
memory[3219] = 32'd6855866;
memory[3220] = 32'd2638020;
memory[3221] = 32'd6363501;
memory[3222] = 32'd7758874;
memory[3223] = 32'd6423611;
memory[3224] = 32'd4483445;
memory[3225] = 32'd6220943;
memory[3226] = 32'd644815;
memory[3227] = 32'd3598167;
memory[3228] = 32'd1539847;
memory[3229] = 32'd691643;
memory[3230] = 32'd7964193;
memory[3231] = 32'd1572322;
memory[3232] = 32'd9076780;
memory[3233] = 32'd2852617;
memory[3234] = 32'd5119204;
memory[3235] = 32'd214107;
memory[3236] = 32'd4460396;
memory[3237] = 32'd8756298;
memory[3238] = 32'd1361591;
memory[3239] = 32'd6416008;
memory[3240] = 32'd6162289;
memory[3241] = 32'd7085193;
memory[3242] = 32'd2833817;
memory[3243] = 32'd6410762;
memory[3244] = 32'd4617267;
memory[3245] = 32'd2795150;
memory[3246] = 32'd4730116;
memory[3247] = 32'd2723354;
memory[3248] = 32'd6270887;
memory[3249] = 32'd9306240;
memory[3250] = 32'd2095572;
memory[3251] = 32'd1425259;
memory[3252] = 32'd5669741;
memory[3253] = 32'd9854446;
memory[3254] = 32'd365223;
memory[3255] = 32'd2669538;
memory[3256] = 32'd8591742;
memory[3257] = 32'd1010038;
memory[3258] = 32'd6267705;
memory[3259] = 32'd131589;
memory[3260] = 32'd1701682;
memory[3261] = 32'd6748250;
memory[3262] = 32'd4220263;
memory[3263] = 32'd3294814;
memory[3264] = 32'd9600867;
memory[3265] = 32'd9339467;
memory[3266] = 32'd3508921;
memory[3267] = 32'd6577616;
memory[3268] = 32'd8095765;
memory[3269] = 32'd7386865;
memory[3270] = 32'd2993624;
memory[3271] = 32'd6774406;
memory[3272] = 32'd4472058;
memory[3273] = 32'd5827441;
memory[3274] = 32'd5701520;
memory[3275] = 32'd9089325;
memory[3276] = 32'd8622591;
memory[3277] = 32'd2947988;
memory[3278] = 32'd1812679;
memory[3279] = 32'd7409831;
memory[3280] = 32'd2254228;
memory[3281] = 32'd3908251;
memory[3282] = 32'd8835090;
memory[3283] = 32'd7923969;
memory[3284] = 32'd3762697;
memory[3285] = 32'd9200313;
memory[3286] = 32'd3109859;
memory[3287] = 32'd4870791;
memory[3288] = 32'd210352;
memory[3289] = 32'd1893916;
memory[3290] = 32'd7518732;
memory[3291] = 32'd4428386;
memory[3292] = 32'd8642166;
memory[3293] = 32'd1738995;
memory[3294] = 32'd7723200;
memory[3295] = 32'd759385;
memory[3296] = 32'd3594814;
memory[3297] = 32'd3748473;
memory[3298] = 32'd7337001;
memory[3299] = 32'd1690579;
memory[3300] = 32'd1135338;
memory[3301] = 32'd2846977;
memory[3302] = 32'd981337;
memory[3303] = 32'd5607396;
memory[3304] = 32'd8674418;
memory[3305] = 32'd6682857;
memory[3306] = 32'd7213073;
memory[3307] = 32'd9813362;
memory[3308] = 32'd9630845;
memory[3309] = 32'd1542104;
memory[3310] = 32'd7223193;
memory[3311] = 32'd4401425;
memory[3312] = 32'd7966707;
memory[3313] = 32'd8574635;
memory[3314] = 32'd4841746;
memory[3315] = 32'd1729405;
memory[3316] = 32'd7774949;
memory[3317] = 32'd7951605;
memory[3318] = 32'd9116548;
memory[3319] = 32'd501653;
memory[3320] = 32'd2361873;
memory[3321] = 32'd6635281;
memory[3322] = 32'd4930039;
memory[3323] = 32'd1004039;
memory[3324] = 32'd8374276;
memory[3325] = 32'd5169591;
memory[3326] = 32'd4279777;
memory[3327] = 32'd1969091;
memory[3328] = 32'd8918064;
memory[3329] = 32'd4133130;
memory[3330] = 32'd6176022;
memory[3331] = 32'd2569755;
memory[3332] = 32'd6980108;
memory[3333] = 32'd7157360;
memory[3334] = 32'd8177151;
memory[3335] = 32'd5654526;
memory[3336] = 32'd6356569;
memory[3337] = 32'd7906577;
memory[3338] = 32'd7984240;
memory[3339] = 32'd5987415;
memory[3340] = 32'd9448681;
memory[3341] = 32'd5207433;
memory[3342] = 32'd2905192;
memory[3343] = 32'd7415389;
memory[3344] = 32'd3782069;
memory[3345] = 32'd7746939;
memory[3346] = 32'd1661146;
memory[3347] = 32'd4073370;
memory[3348] = 32'd8214896;
memory[3349] = 32'd777694;
memory[3350] = 32'd4575023;
memory[3351] = 32'd576770;
memory[3352] = 32'd7412975;
memory[3353] = 32'd2021414;
memory[3354] = 32'd4097161;
memory[3355] = 32'd8303604;
memory[3356] = 32'd7191005;
memory[3357] = 32'd8376938;
memory[3358] = 32'd272695;
memory[3359] = 32'd8625421;
memory[3360] = 32'd2510069;
memory[3361] = 32'd8965069;
memory[3362] = 32'd1195176;
memory[3363] = 32'd9490177;
memory[3364] = 32'd6122429;
memory[3365] = 32'd1888680;
memory[3366] = 32'd7661055;
memory[3367] = 32'd2478999;
memory[3368] = 32'd9795257;
memory[3369] = 32'd5645296;
memory[3370] = 32'd982766;
memory[3371] = 32'd9243938;
memory[3372] = 32'd3369081;
memory[3373] = 32'd3887958;
memory[3374] = 32'd9175679;
memory[3375] = 32'd9667502;
memory[3376] = 32'd4151249;
memory[3377] = 32'd836825;
memory[3378] = 32'd6257224;
memory[3379] = 32'd2366146;
memory[3380] = 32'd4130872;
memory[3381] = 32'd832247;
memory[3382] = 32'd2942916;
memory[3383] = 32'd1543847;
memory[3384] = 32'd2853661;
memory[3385] = 32'd7040077;
memory[3386] = 32'd9847451;
memory[3387] = 32'd2561018;
memory[3388] = 32'd5417016;
memory[3389] = 32'd2636498;
memory[3390] = 32'd1186440;
memory[3391] = 32'd443437;
memory[3392] = 32'd1601568;
memory[3393] = 32'd2381616;
memory[3394] = 32'd2449966;
memory[3395] = 32'd240349;
memory[3396] = 32'd4270296;
memory[3397] = 32'd111021;
memory[3398] = 32'd2719348;
memory[3399] = 32'd6581905;
memory[3400] = 32'd8272669;
memory[3401] = 32'd6218466;
memory[3402] = 32'd8342196;
memory[3403] = 32'd1641751;
memory[3404] = 32'd2622777;
memory[3405] = 32'd7517875;
memory[3406] = 32'd3825605;
memory[3407] = 32'd6774026;
memory[3408] = 32'd871053;
memory[3409] = 32'd82830;
memory[3410] = 32'd9140172;
memory[3411] = 32'd5001925;
memory[3412] = 32'd3431429;
memory[3413] = 32'd2083088;
memory[3414] = 32'd6545772;
memory[3415] = 32'd8801443;
memory[3416] = 32'd1639518;
memory[3417] = 32'd8909576;
memory[3418] = 32'd1362461;
memory[3419] = 32'd9572886;
memory[3420] = 32'd4062426;
memory[3421] = 32'd2548901;
memory[3422] = 32'd16323;
memory[3423] = 32'd5663994;
memory[3424] = 32'd7446870;
memory[3425] = 32'd2466289;
memory[3426] = 32'd8420696;
memory[3427] = 32'd4233518;
memory[3428] = 32'd5093662;
memory[3429] = 32'd3656396;
memory[3430] = 32'd815424;
memory[3431] = 32'd3366332;
memory[3432] = 32'd9874863;
memory[3433] = 32'd9157620;
memory[3434] = 32'd7524435;
memory[3435] = 32'd2497640;
memory[3436] = 32'd9191847;
memory[3437] = 32'd3866392;
memory[3438] = 32'd1788018;
memory[3439] = 32'd62900;
memory[3440] = 32'd3949222;
memory[3441] = 32'd3444543;
memory[3442] = 32'd5064825;
memory[3443] = 32'd9897004;
memory[3444] = 32'd8043983;
memory[3445] = 32'd4126950;
memory[3446] = 32'd8698447;
memory[3447] = 32'd9683501;
memory[3448] = 32'd5552878;
memory[3449] = 32'd60908;
memory[3450] = 32'd9256387;
memory[3451] = 32'd9615304;
memory[3452] = 32'd5126162;
memory[3453] = 32'd1789062;
memory[3454] = 32'd7795651;
memory[3455] = 32'd2573032;
memory[3456] = 32'd4255351;
memory[3457] = 32'd6216347;
memory[3458] = 32'd9322902;
memory[3459] = 32'd1865366;
memory[3460] = 32'd9872743;
memory[3461] = 32'd138326;
memory[3462] = 32'd7748050;
memory[3463] = 32'd2263958;
memory[3464] = 32'd1812298;
memory[3465] = 32'd7788837;
memory[3466] = 32'd7277950;
memory[3467] = 32'd3520498;
memory[3468] = 32'd1655229;
memory[3469] = 32'd9065969;
memory[3470] = 32'd3583398;
memory[3471] = 32'd8120804;
memory[3472] = 32'd2510512;
memory[3473] = 32'd1164576;
memory[3474] = 32'd8017808;
memory[3475] = 32'd3070847;
memory[3476] = 32'd7807878;
memory[3477] = 32'd6716255;
memory[3478] = 32'd2754349;
memory[3479] = 32'd5877108;
memory[3480] = 32'd6777163;
memory[3481] = 32'd2010736;
memory[3482] = 32'd8008764;
memory[3483] = 32'd4419677;
memory[3484] = 32'd6316151;
memory[3485] = 32'd5804415;
memory[3486] = 32'd6992709;
memory[3487] = 32'd3087854;
memory[3488] = 32'd4537114;
memory[3489] = 32'd6315612;
memory[3490] = 32'd4953220;
memory[3491] = 32'd6926210;
memory[3492] = 32'd8970290;
memory[3493] = 32'd2701270;
memory[3494] = 32'd9190168;
memory[3495] = 32'd3298941;
memory[3496] = 32'd490107;
memory[3497] = 32'd8984471;
memory[3498] = 32'd6819439;
memory[3499] = 32'd4661689;
memory[3500] = 32'd8050440;
memory[3501] = 32'd2919189;
memory[3502] = 32'd2782493;
memory[3503] = 32'd3077304;
memory[3504] = 32'd6600117;
memory[3505] = 32'd3316653;
memory[3506] = 32'd6148151;
memory[3507] = 32'd6924347;
memory[3508] = 32'd32908;
memory[3509] = 32'd1418852;
memory[3510] = 32'd2801455;
memory[3511] = 32'd9326423;
memory[3512] = 32'd5945941;
memory[3513] = 32'd3326572;
memory[3514] = 32'd3746101;
memory[3515] = 32'd2262092;
memory[3516] = 32'd1647339;
memory[3517] = 32'd3255162;
memory[3518] = 32'd5349946;
memory[3519] = 32'd6184454;
memory[3520] = 32'd2087126;
memory[3521] = 32'd2819519;
memory[3522] = 32'd5627016;
memory[3523] = 32'd3573769;
memory[3524] = 32'd5520789;
memory[3525] = 32'd4817184;
memory[3526] = 32'd6872710;
memory[3527] = 32'd8527249;
memory[3528] = 32'd3801655;
memory[3529] = 32'd6208501;
memory[3530] = 32'd5705290;
memory[3531] = 32'd4368447;
memory[3532] = 32'd1644042;
memory[3533] = 32'd8487783;
memory[3534] = 32'd9962103;
memory[3535] = 32'd760512;
memory[3536] = 32'd4320788;
memory[3537] = 32'd8626607;
memory[3538] = 32'd201211;
memory[3539] = 32'd4353696;
memory[3540] = 32'd2561811;
memory[3541] = 32'd5519019;
memory[3542] = 32'd6196471;
memory[3543] = 32'd8507752;
memory[3544] = 32'd8845591;
memory[3545] = 32'd2458924;
memory[3546] = 32'd3286196;
memory[3547] = 32'd492930;
memory[3548] = 32'd5714087;
memory[3549] = 32'd8636143;
memory[3550] = 32'd9193736;
memory[3551] = 32'd317565;
memory[3552] = 32'd1455662;
memory[3553] = 32'd4820752;
memory[3554] = 32'd3891334;
memory[3555] = 32'd9492803;
memory[3556] = 32'd2154289;
memory[3557] = 32'd3280396;
memory[3558] = 32'd536404;
memory[3559] = 32'd8472296;
memory[3560] = 32'd9488897;
memory[3561] = 32'd6241694;
memory[3562] = 32'd5357096;
memory[3563] = 32'd3649292;
memory[3564] = 32'd7245829;
memory[3565] = 32'd5319199;
memory[3566] = 32'd6926156;
memory[3567] = 32'd1566617;
memory[3568] = 32'd6462158;
memory[3569] = 32'd7127367;
memory[3570] = 32'd8436665;
memory[3571] = 32'd1540322;
memory[3572] = 32'd2646386;
memory[3573] = 32'd4633137;
memory[3574] = 32'd48074;
memory[3575] = 32'd1491977;
memory[3576] = 32'd7092061;
memory[3577] = 32'd3334271;
memory[3578] = 32'd1984908;
memory[3579] = 32'd5322500;
memory[3580] = 32'd4486766;
memory[3581] = 32'd3694996;
memory[3582] = 32'd5640066;
memory[3583] = 32'd8458780;
memory[3584] = 32'd8515749;
memory[3585] = 32'd9531400;
memory[3586] = 32'd467935;
memory[3587] = 32'd670038;
memory[3588] = 32'd2811797;
memory[3589] = 32'd1004340;
memory[3590] = 32'd9142334;
memory[3591] = 32'd4817046;
memory[3592] = 32'd9762386;
memory[3593] = 32'd4499430;
memory[3594] = 32'd982690;
memory[3595] = 32'd7008216;
memory[3596] = 32'd2334982;
memory[3597] = 32'd7908846;
memory[3598] = 32'd1091185;
memory[3599] = 32'd1313492;
memory[3600] = 32'd5036214;
memory[3601] = 32'd9527851;
memory[3602] = 32'd2853814;
memory[3603] = 32'd198952;
memory[3604] = 32'd6677340;
memory[3605] = 32'd5418241;
memory[3606] = 32'd1690930;
memory[3607] = 32'd6285753;
memory[3608] = 32'd1268864;
memory[3609] = 32'd6192190;
memory[3610] = 32'd1608254;
memory[3611] = 32'd5755630;
memory[3612] = 32'd9887186;
memory[3613] = 32'd9764672;
memory[3614] = 32'd6730762;
memory[3615] = 32'd919287;
memory[3616] = 32'd9296072;
memory[3617] = 32'd7198697;
memory[3618] = 32'd1589325;
memory[3619] = 32'd4624221;
memory[3620] = 32'd719389;
memory[3621] = 32'd731660;
memory[3622] = 32'd1957620;
memory[3623] = 32'd481776;
memory[3624] = 32'd7747442;
memory[3625] = 32'd2940310;
memory[3626] = 32'd7489992;
memory[3627] = 32'd82424;
memory[3628] = 32'd3365509;
memory[3629] = 32'd1097529;
memory[3630] = 32'd3912269;
memory[3631] = 32'd918075;
memory[3632] = 32'd625380;
memory[3633] = 32'd6766083;
memory[3634] = 32'd1117027;
memory[3635] = 32'd7302720;
memory[3636] = 32'd2184324;
memory[3637] = 32'd5324309;
memory[3638] = 32'd3588474;
memory[3639] = 32'd3453188;
memory[3640] = 32'd1516499;
memory[3641] = 32'd7713080;
memory[3642] = 32'd1725170;
memory[3643] = 32'd3920038;
memory[3644] = 32'd7477752;
memory[3645] = 32'd8455932;
memory[3646] = 32'd4839325;
memory[3647] = 32'd9290176;
memory[3648] = 32'd8170982;
memory[3649] = 32'd6428651;
memory[3650] = 32'd3914398;
memory[3651] = 32'd8890371;
memory[3652] = 32'd9676663;
memory[3653] = 32'd8388370;
memory[3654] = 32'd9372147;
memory[3655] = 32'd9940457;
memory[3656] = 32'd3845032;
memory[3657] = 32'd9378491;
memory[3658] = 32'd2539234;
memory[3659] = 32'd7210541;
memory[3660] = 32'd476021;
memory[3661] = 32'd6451503;
memory[3662] = 32'd8128616;
memory[3663] = 32'd3617753;
memory[3664] = 32'd5733938;
memory[3665] = 32'd1761996;
memory[3666] = 32'd3436826;
memory[3667] = 32'd7918263;
memory[3668] = 32'd7086305;
memory[3669] = 32'd9541652;
memory[3670] = 32'd3887803;
memory[3671] = 32'd1119157;
memory[3672] = 32'd7254732;
memory[3673] = 32'd8129326;
memory[3674] = 32'd5039195;
memory[3675] = 32'd7248836;
memory[3676] = 32'd6585258;
memory[3677] = 32'd9878520;
memory[3678] = 32'd6539012;
memory[3679] = 32'd7272592;
memory[3680] = 32'd8823523;
memory[3681] = 32'd2969762;
memory[3682] = 32'd6162964;
memory[3683] = 32'd1016538;
memory[3684] = 32'd1358132;
memory[3685] = 32'd8051463;
memory[3686] = 32'd3473348;
memory[3687] = 32'd5203165;
memory[3688] = 32'd9946307;
memory[3689] = 32'd6012582;
memory[3690] = 32'd4930058;
memory[3691] = 32'd422328;
memory[3692] = 32'd4980437;
memory[3693] = 32'd5575027;
memory[3694] = 32'd6556433;
memory[3695] = 32'd714375;
memory[3696] = 32'd7337023;
memory[3697] = 32'd9993259;
memory[3698] = 32'd1148990;
memory[3699] = 32'd4423328;
memory[3700] = 32'd9534911;
memory[3701] = 32'd7553146;
memory[3702] = 32'd5542485;
memory[3703] = 32'd9305995;
memory[3704] = 32'd5682472;
memory[3705] = 32'd3098032;
memory[3706] = 32'd6554831;
memory[3707] = 32'd4784082;
memory[3708] = 32'd5492905;
memory[3709] = 32'd5610196;
memory[3710] = 32'd2056675;
memory[3711] = 32'd4316428;
memory[3712] = 32'd8579958;
memory[3713] = 32'd8219639;
memory[3714] = 32'd7849319;
memory[3715] = 32'd2454443;
memory[3716] = 32'd8787454;
memory[3717] = 32'd1322667;
memory[3718] = 32'd173960;
memory[3719] = 32'd8733761;
memory[3720] = 32'd9851601;
memory[3721] = 32'd7620370;
memory[3722] = 32'd1672441;
memory[3723] = 32'd4832038;
memory[3724] = 32'd3195397;
memory[3725] = 32'd8228875;
memory[3726] = 32'd5546413;
memory[3727] = 32'd532420;
memory[3728] = 32'd738486;
memory[3729] = 32'd9211756;
memory[3730] = 32'd7472101;
memory[3731] = 32'd273398;
memory[3732] = 32'd6764902;
memory[3733] = 32'd5530938;
memory[3734] = 32'd2095745;
memory[3735] = 32'd2447374;
memory[3736] = 32'd1145323;
memory[3737] = 32'd1166929;
memory[3738] = 32'd7231456;
memory[3739] = 32'd6638228;
memory[3740] = 32'd6777125;
memory[3741] = 32'd9288131;
memory[3742] = 32'd3471008;
memory[3743] = 32'd7873435;
memory[3744] = 32'd24122;
memory[3745] = 32'd3836679;
memory[3746] = 32'd2844230;
memory[3747] = 32'd8811577;
memory[3748] = 32'd5159346;
memory[3749] = 32'd3018190;
memory[3750] = 32'd61690;
memory[3751] = 32'd5010947;
memory[3752] = 32'd3154913;
memory[3753] = 32'd1734132;
memory[3754] = 32'd2359337;
memory[3755] = 32'd6350310;
memory[3756] = 32'd9963007;
memory[3757] = 32'd7905751;
memory[3758] = 32'd9399083;
memory[3759] = 32'd701493;
memory[3760] = 32'd7117507;
memory[3761] = 32'd9387536;
memory[3762] = 32'd3491243;
memory[3763] = 32'd3882409;
memory[3764] = 32'd7434826;
memory[3765] = 32'd5586989;
memory[3766] = 32'd8846135;
memory[3767] = 32'd8580149;
memory[3768] = 32'd6753918;
memory[3769] = 32'd6077591;
memory[3770] = 32'd5218377;
memory[3771] = 32'd6047395;
memory[3772] = 32'd5365723;
memory[3773] = 32'd1205738;
memory[3774] = 32'd3920830;
memory[3775] = 32'd7906197;
memory[3776] = 32'd5042417;
memory[3777] = 32'd9281413;
memory[3778] = 32'd6717774;
memory[3779] = 32'd2718116;
memory[3780] = 32'd4815955;
memory[3781] = 32'd6779465;
memory[3782] = 32'd245415;
memory[3783] = 32'd7970868;
memory[3784] = 32'd1029949;
memory[3785] = 32'd2604753;
memory[3786] = 32'd4321179;
memory[3787] = 32'd992956;
memory[3788] = 32'd3026856;
memory[3789] = 32'd6236614;
memory[3790] = 32'd4210801;
memory[3791] = 32'd2660715;
memory[3792] = 32'd5624150;
memory[3793] = 32'd218397;
memory[3794] = 32'd9059476;
memory[3795] = 32'd3058976;
memory[3796] = 32'd8321738;
memory[3797] = 32'd7905611;
memory[3798] = 32'd1639126;
memory[3799] = 32'd7592008;
memory[3800] = 32'd3983202;
memory[3801] = 32'd9373855;
memory[3802] = 32'd3639403;
memory[3803] = 32'd1865277;
memory[3804] = 32'd579593;
memory[3805] = 32'd76585;
memory[3806] = 32'd9771475;
memory[3807] = 32'd5622011;
memory[3808] = 32'd9357998;
memory[3809] = 32'd9005601;
memory[3810] = 32'd8340127;
memory[3811] = 32'd6690306;
memory[3812] = 32'd8301418;
memory[3813] = 32'd8585542;
memory[3814] = 32'd4661174;
memory[3815] = 32'd9331367;
memory[3816] = 32'd3706647;
memory[3817] = 32'd8982353;
memory[3818] = 32'd324323;
memory[3819] = 32'd6733503;
memory[3820] = 32'd5218967;
memory[3821] = 32'd7051477;
memory[3822] = 32'd9394218;
memory[3823] = 32'd3359469;
memory[3824] = 32'd9786226;
memory[3825] = 32'd8453694;
memory[3826] = 32'd6418446;
memory[3827] = 32'd8107964;
memory[3828] = 32'd6359305;
memory[3829] = 32'd573924;
memory[3830] = 32'd5699972;
memory[3831] = 32'd2858860;
memory[3832] = 32'd9947779;
memory[3833] = 32'd1855727;
memory[3834] = 32'd4724137;
memory[3835] = 32'd3043725;
memory[3836] = 32'd4448664;
memory[3837] = 32'd7011964;
memory[3838] = 32'd8665736;
memory[3839] = 32'd6323015;
memory[3840] = 32'd6017566;
memory[3841] = 32'd9522215;
memory[3842] = 32'd3013321;
memory[3843] = 32'd4318984;
memory[3844] = 32'd624109;
memory[3845] = 32'd7674495;
memory[3846] = 32'd3650352;
memory[3847] = 32'd4330757;
memory[3848] = 32'd9173201;
memory[3849] = 32'd6491027;
memory[3850] = 32'd1064260;
memory[3851] = 32'd6908520;
memory[3852] = 32'd6058856;
memory[3853] = 32'd2974831;
memory[3854] = 32'd267990;
memory[3855] = 32'd5845082;
memory[3856] = 32'd1428525;
memory[3857] = 32'd9202788;
memory[3858] = 32'd3953046;
memory[3859] = 32'd304183;
memory[3860] = 32'd9776712;
memory[3861] = 32'd2169370;
memory[3862] = 32'd3163043;
memory[3863] = 32'd9724491;
memory[3864] = 32'd6541449;
memory[3865] = 32'd403532;
memory[3866] = 32'd2768216;
memory[3867] = 32'd3506466;
memory[3868] = 32'd7415497;
memory[3869] = 32'd3950304;
memory[3870] = 32'd9829481;
memory[3871] = 32'd3433063;
memory[3872] = 32'd5988871;
memory[3873] = 32'd5359154;
memory[3874] = 32'd268399;
memory[3875] = 32'd6612981;
memory[3876] = 32'd5550001;
memory[3877] = 32'd3918751;
memory[3878] = 32'd3460090;
memory[3879] = 32'd4723202;
memory[3880] = 32'd2926131;
memory[3881] = 32'd7040702;
memory[3882] = 32'd4148075;
memory[3883] = 32'd8984987;
memory[3884] = 32'd15533;
memory[3885] = 32'd4416065;
memory[3886] = 32'd4830070;
memory[3887] = 32'd3960411;
memory[3888] = 32'd6135205;
memory[3889] = 32'd1299468;
memory[3890] = 32'd6780946;
memory[3891] = 32'd5911917;
memory[3892] = 32'd5985191;
memory[3893] = 32'd9943989;
memory[3894] = 32'd8152760;
memory[3895] = 32'd5042992;
memory[3896] = 32'd2863873;
memory[3897] = 32'd3437329;
memory[3898] = 32'd8549458;
memory[3899] = 32'd279370;
memory[3900] = 32'd7387633;
memory[3901] = 32'd895291;
memory[3902] = 32'd6228785;
memory[3903] = 32'd5892857;
memory[3904] = 32'd8770797;
memory[3905] = 32'd9013537;
memory[3906] = 32'd5022190;
memory[3907] = 32'd4320799;
memory[3908] = 32'd2932288;
memory[3909] = 32'd8482280;
memory[3910] = 32'd1560353;
memory[3911] = 32'd8374771;
memory[3912] = 32'd8039334;
memory[3913] = 32'd5708428;
memory[3914] = 32'd7359759;
memory[3915] = 32'd571220;
memory[3916] = 32'd2640845;
memory[3917] = 32'd4706181;
memory[3918] = 32'd7047983;
memory[3919] = 32'd8776050;
memory[3920] = 32'd8522001;
memory[3921] = 32'd3828929;
memory[3922] = 32'd7204319;
memory[3923] = 32'd4507192;
memory[3924] = 32'd6289270;
memory[3925] = 32'd5357080;
memory[3926] = 32'd2066537;
memory[3927] = 32'd9153143;
memory[3928] = 32'd8794409;
memory[3929] = 32'd3132347;
memory[3930] = 32'd1948866;
memory[3931] = 32'd8698394;
memory[3932] = 32'd4027639;
memory[3933] = 32'd694003;
memory[3934] = 32'd7107603;
memory[3935] = 32'd5314788;
memory[3936] = 32'd9707540;
memory[3937] = 32'd2129793;
memory[3938] = 32'd9635587;
memory[3939] = 32'd5156181;
memory[3940] = 32'd3128425;
memory[3941] = 32'd1195941;
memory[3942] = 32'd3530952;
memory[3943] = 32'd3684112;
memory[3944] = 32'd9420721;
memory[3945] = 32'd3407063;
memory[3946] = 32'd4255332;
memory[3947] = 32'd2061567;
memory[3948] = 32'd8113244;
memory[3949] = 32'd1303315;
memory[3950] = 32'd3353969;
memory[3951] = 32'd6635246;
memory[3952] = 32'd5132244;
memory[3953] = 32'd558289;
memory[3954] = 32'd3658790;
memory[3955] = 32'd1421514;
memory[3956] = 32'd8431721;
memory[3957] = 32'd5725327;
memory[3958] = 32'd3091009;
memory[3959] = 32'd7226130;
memory[3960] = 32'd8857675;
memory[3961] = 32'd5039875;
memory[3962] = 32'd8440876;
memory[3963] = 32'd5401666;
memory[3964] = 32'd8250231;
memory[3965] = 32'd5548480;
memory[3966] = 32'd716454;
memory[3967] = 32'd7957771;
memory[3968] = 32'd194625;
memory[3969] = 32'd352042;
memory[3970] = 32'd5630304;
memory[3971] = 32'd5839403;
memory[3972] = 32'd4064335;
memory[3973] = 32'd9161257;
memory[3974] = 32'd9523515;
memory[3975] = 32'd3485056;
memory[3976] = 32'd5084672;
memory[3977] = 32'd3778847;
memory[3978] = 32'd8062975;
memory[3979] = 32'd3197917;
memory[3980] = 32'd7598514;
memory[3981] = 32'd1416945;
memory[3982] = 32'd9833163;
memory[3983] = 32'd2730758;
memory[3984] = 32'd4491586;
memory[3985] = 32'd3491953;
memory[3986] = 32'd6668624;
memory[3987] = 32'd2923307;
memory[3988] = 32'd9217281;
memory[3989] = 32'd9759633;
memory[3990] = 32'd2665789;
memory[3991] = 32'd591308;
memory[3992] = 32'd7315861;
memory[3993] = 32'd3623017;
memory[3994] = 32'd5992974;
memory[3995] = 32'd5566092;
memory[3996] = 32'd1687849;
memory[3997] = 32'd6709428;
memory[3998] = 32'd6040215;
memory[3999] = 32'd1882475;
memory[4000] = 32'd9577822;
memory[4001] = 32'd4186872;
memory[4002] = 32'd238230;
memory[4003] = 32'd3642157;
memory[4004] = 32'd5864481;
memory[4005] = 32'd9761745;
memory[4006] = 32'd9643566;
memory[4007] = 32'd949153;
memory[4008] = 32'd3540592;
memory[4009] = 32'd7706541;
memory[4010] = 32'd4147070;
memory[4011] = 32'd3655458;
memory[4012] = 32'd1639838;
memory[4013] = 32'd6496585;
memory[4014] = 32'd6386216;
memory[4015] = 32'd6131424;
memory[4016] = 32'd9988539;
memory[4017] = 32'd5571192;
memory[4018] = 32'd1571083;
memory[4019] = 32'd1722172;
memory[4020] = 32'd7847177;
memory[4021] = 32'd4236872;
memory[4022] = 32'd4829832;
memory[4023] = 32'd5163038;
memory[4024] = 32'd376242;
memory[4025] = 32'd822806;
memory[4026] = 32'd3245482;
memory[4027] = 32'd2064091;
memory[4028] = 32'd48586;
memory[4029] = 32'd1802050;
memory[4030] = 32'd6462918;
memory[4031] = 32'd9626409;
memory[4032] = 32'd5988922;
memory[4033] = 32'd6701148;
memory[4034] = 32'd5784918;
memory[4035] = 32'd4369755;
memory[4036] = 32'd8979245;
memory[4037] = 32'd5428484;
memory[4038] = 32'd5318908;
memory[4039] = 32'd5036189;
memory[4040] = 32'd5651378;
memory[4041] = 32'd9465979;
memory[4042] = 32'd8691647;
memory[4043] = 32'd7291216;
memory[4044] = 32'd5962564;
memory[4045] = 32'd7594215;
memory[4046] = 32'd5938993;
memory[4047] = 32'd8467455;
memory[4048] = 32'd3165407;
memory[4049] = 32'd7510076;
memory[4050] = 32'd2705979;
memory[4051] = 32'd1012585;
memory[4052] = 32'd4263301;
memory[4053] = 32'd7535811;
memory[4054] = 32'd8691975;
memory[4055] = 32'd7155895;
memory[4056] = 32'd874969;
memory[4057] = 32'd4453810;
memory[4058] = 32'd9219986;
memory[4059] = 32'd923556;
memory[4060] = 32'd8772212;
memory[4061] = 32'd8199257;
memory[4062] = 32'd3066317;
memory[4063] = 32'd7277486;
memory[4064] = 32'd7416757;
memory[4065] = 32'd8851235;
memory[4066] = 32'd1647241;
memory[4067] = 32'd6396003;
memory[4068] = 32'd6796072;
memory[4069] = 32'd6966149;
memory[4070] = 32'd1432192;
memory[4071] = 32'd2447450;
memory[4072] = 32'd8948480;
memory[4073] = 32'd123840;
memory[4074] = 32'd2255018;
memory[4075] = 32'd7427397;
memory[4076] = 32'd7718055;
memory[4077] = 32'd8194011;
memory[4078] = 32'd8411204;
memory[4079] = 32'd3399815;
memory[4080] = 32'd8220440;
memory[4081] = 32'd1117184;
memory[4082] = 32'd4412400;
memory[4083] = 32'd5000093;
memory[4084] = 32'd1169347;
memory[4085] = 32'd5620727;
memory[4086] = 32'd2155988;
memory[4087] = 32'd2044317;
memory[4088] = 32'd74537;
memory[4089] = 32'd1375974;
memory[4090] = 32'd2967873;
memory[4091] = 32'd1363101;
memory[4092] = 32'd2091583;
memory[4093] = 32'd6034190;
memory[4094] = 32'd8640587;
memory[4095] = 32'd9508341;

end

endmodule
